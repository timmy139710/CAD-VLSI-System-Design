// Verilog HDL NetList 
//   timeStamp 2005 7 28 16 6 31 
//   author "Avanti Corporation."
//   program "A2Hdl" 
//   design library: io_tpd013n3
//   cell name     : io_tpd013n3.CEL (version 1)
module PVDD1CDG ();
endmodule 
module PVDD2CDG ();
endmodule 
module PVDD2POC ();
endmodule 
module PVSS1CDG ();
endmodule 
module PVSS2CDG ();
endmodule 
module PVSS3CDG ();
endmodule 
module PXOE1CDG ( XC , XE , XI , XO );
    output XC ;
    input XE ;
    input XI ;
    output XO ;
endmodule 
module PXOE2CDG ( XC , XE , XI , XO );
    output XC ;
    input XE ;
    input XI ;
    output XO ;
endmodule 
module PAD60N ();
endmodule 
module PCORNERN ();
endmodule 
module PDC0102CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PDC0204CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PDC0408CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PDC1216CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PDS0102CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PDS0204CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PDS0408CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PDS1216CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PFEED0005N ();
endmodule 
module PFEED001N ();
endmodule 
module PFEED01N ();
endmodule 
module PFEED10N ();
endmodule 
module PFEED1N ();
endmodule 
module PFEED20N ();
endmodule 
module PFEED5N ();
endmodule 
module PRC0102CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PRC0204CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PRC0408CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PRC1216CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PRS0102CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PRS0204CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PRS0408CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 
module PRS1216CDG ( C , DS , I , IE , OEN , PAD , PE , PS );
    output C ;
    input DS ;
    input I ;
    input IE ;
    input OEN ;
    inout PAD ;
    input PE ;
    input PS ;
endmodule 

