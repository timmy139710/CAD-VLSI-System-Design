.SUBCKT RF2SH64x16
+ QA[0] QA[1] QA[2] QA[3] QA[4] QA[5] QA[6] QA[7] QA[8] QA[9] QA[10] QA[11] QA[12] QA[13] QA[14] QA[15] 
+ CLKA CENA 
+ AA[0] AA[1] AA[2] AA[3] AA[4] AA[5]
+ AB[0] AB[1] AB[2] AB[3] AB[4] AB[5] 
+ DB[0] DB[1] DB[2] DB[3] DB[4] DB[5] DB[6] DB[7] DB[8] DB[9] DB[10] DB[11] DB[12] DB[13] DB[14] DB[15] 
+ CLKB CENB 
+ VDD VSS
.ENDS
