// Verilog HDL NetList 
//   timeStamp 2005 7 28 16 16 54 
//   author "Avanti Corporation."
//   program "A2Hdl" 
//   design library: io_tpz013g3
//   cell name     : io_tpz013g3.CEL (version 1)
module PDUWDGZ ( C , PAD , REN );
    output C ;
    input PAD ;
    input REN ;
endmodule 
module PDXO01DG ( XC , XIN , XOUT );
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDXO02DG ( XC , XIN , XOUT );
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDXO03DG ( XC , XIN , XOUT );
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDXOE1DG ( E , XC , XIN , XOUT );
    input E ;
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDXOE2DG ( E , XC , XIN , XOUT );
    input E ;
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDXOE3DG ( E , XC , XIN , XOUT );
    input E ;
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PFEED0_005Z ();
endmodule 
module PFEED0_01Z ();
endmodule 
module PDD12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDDDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDDSDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDDW02DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW04DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW08DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW12DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW16DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRD24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRDW08DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRDW12DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRDW16DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRDW24DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRO08CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PRO12CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PRO16CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PRO24CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDU02DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU02SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU04DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU04SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDUDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDUSDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDUW02DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW04DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW08DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW12DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW16DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW24DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRUW12DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRUW16DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRUW24DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PVDD1DGZ ();
endmodule 
module PVDD2DGZ ();
endmodule 
module PVDD2POC ();
endmodule 
module PVSS1DGZ ();
endmodule 
module PVSS2DGZ ();
endmodule 
module PVSS3DGZ ();
endmodule 
module PFEED0_1Z ();
endmodule 
module PFEED10Z ();
endmodule 
module PFEED1Z ();
endmodule 
module PFEED20Z ();
endmodule 
module PFEED5Z ();
endmodule 
module PRB08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB04DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB04SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD02DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD02SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD04DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD04SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRT08DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PRT12DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PRT16DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PRT24DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PRU08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRUW08DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW24DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDWDGZ ( C , PAD , REN );
    output C ;
    input PAD ;
    input REN ;
endmodule 
module PDIDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDISDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDO02CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO04CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO08CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO12CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO16CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO24CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDT02DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDT04DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDT08DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDT12DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDT16DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDT24DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PADIZ40 ();
endmodule 
module PADIZ45 ();
endmodule 
module PADLZ60 ();
endmodule 
module PADLZ85 ();
endmodule 
module PADOZ40 ();
endmodule 
module PADOZ45 ();
endmodule 
module PCI33DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PCI33SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PCI66DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PCI66SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PCORNERDGZ ();
endmodule 
module PDB02DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB02SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 

