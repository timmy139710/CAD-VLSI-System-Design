module RF2SH64x16 (
   QA,
   AA,
   CLKA,
   CENA,
   AB,
   DB,
   CLKB,
   CENB
);
   output [15:0] QA;
   input [5:0] AA;
   input CLKA;
   input CENA;
   input [5:0] AB;
   input [15:0] DB;
   input CLKB;
   input CENB;

endmodule
