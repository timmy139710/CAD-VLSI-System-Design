###############################################################################
#TSMC Library/IP Product
#Filename: tpz013g3_8lm.lef
#Technology: CL013G
#Product Type: Standard I/O
#Product Name: tpz013g3
#Version: 210b
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################

###############################################################################
# Modified by CIC 2006/07/05 (CBDK013_TSMC_Artisan v1.1) 
#
# Added METAL1 PIN on PCORNERDGZ Cell for recognizing corner orientation
#
###############################################################################

SITE pad
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 0.005 BY 246.000 ;
END pad 

SITE corner
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 246.000 BY 246.000 ;
END corner

MACRO PADIZ40
    CLASS BLOCK ;
    FOREIGN PADIZ40 17.000 0.000  ;
    ORIGIN -17.000 0.000 ;
    SIZE 35.000 BY 88.800 ;
    SYMMETRY x y r90 ;
    OBS
        LAYER METAL1 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL2 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL3 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL4 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL5 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL6 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL7 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL8 ;
        RECT  17.000 0.000 52.000 88.800 ;
    END
END PADIZ40

MACRO PADIZ45
    CLASS BLOCK ;
    FOREIGN PADIZ45 17.000 0.000  ;
    ORIGIN -17.000 0.000 ;
    SIZE 35.000 BY 88.800 ;
    SYMMETRY x y r90 ;
    OBS
        LAYER METAL1 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL2 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL3 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL4 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL5 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL6 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL7 ;
        RECT  17.000 0.000 52.000 88.800 ;
        LAYER METAL8 ;
        RECT  17.000 0.000 52.000 88.800 ;
    END
END PADIZ45

MACRO PADLZ60
    CLASS BLOCK ;
    FOREIGN PADLZ60 11.000 0.000  ;
    ORIGIN -11.000 0.000 ;
    SIZE 35.000 BY 80.000 ;
    SYMMETRY x y r90 ;
    OBS
        LAYER METAL1 ;
        RECT  11.000 0.000 46.000 80.000 ;
        LAYER METAL2 ;
        RECT  11.000 0.000 46.000 80.000 ;
        LAYER METAL3 ;
        RECT  11.000 0.000 46.000 80.000 ;
        LAYER METAL4 ;
        RECT  11.000 0.000 46.000 80.000 ;
        LAYER METAL5 ;
        RECT  11.000 0.000 46.000 80.000 ;
        LAYER METAL6 ;
        RECT  11.000 0.000 46.000 80.000 ;
        LAYER METAL7 ;
        RECT  11.000 0.000 46.000 80.000 ;
        LAYER METAL8 ;
        RECT  11.000 0.000 46.000 80.000 ;
    END
END PADLZ60

MACRO PADLZ85
    CLASS BLOCK ;
    FOREIGN PADLZ85 22.000 0.000  ;
    ORIGIN -22.000 0.000 ;
    SIZE 35.000 BY 89.000 ;
    SYMMETRY x y r90 ;
    OBS
        LAYER METAL1 ;
        RECT  22.000 0.000 57.000 89.000 ;
        LAYER METAL2 ;
        RECT  22.000 0.000 57.000 89.000 ;
        LAYER METAL3 ;
        RECT  22.000 0.000 57.000 89.000 ;
        LAYER METAL4 ;
        RECT  22.000 0.000 57.000 89.000 ;
        LAYER METAL5 ;
        RECT  22.000 0.000 57.000 89.000 ;
        LAYER METAL6 ;
        RECT  22.000 0.000 57.000 89.000 ;
        LAYER METAL7 ;
        RECT  22.000 0.000 57.000 89.000 ;
        LAYER METAL8 ;
        RECT  22.000 0.000 57.000 89.000 ;
    END
END PADLZ85

MACRO PADOZ40
    CLASS BLOCK ;
    FOREIGN PADOZ40 17.000 0.000  ;
    ORIGIN -17.000 0.000 ;
    SIZE 35.000 BY 203.800 ;
    SYMMETRY x y r90 ;
    OBS
        LAYER METAL1 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL2 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL3 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL4 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL5 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL6 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL7 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL8 ;
        RECT  17.000 0.000 52.000 203.800 ;
    END
END PADOZ40

MACRO PADOZ45
    CLASS BLOCK ;
    FOREIGN PADOZ45 17.000 0.000  ;
    ORIGIN -17.000 0.000 ;
    SIZE 35.000 BY 203.800 ;
    SYMMETRY x y r90 ;
    OBS
        LAYER METAL1 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL2 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL3 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL4 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL5 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL6 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL7 ;
        RECT  17.000 0.000 52.000 203.800 ;
        LAYER METAL8 ;
        RECT  17.000 0.000 52.000 203.800 ;
    END
END PADOZ45

MACRO PCI33DGZ
    CLASS PAD ;
    FOREIGN PCI33DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PCI33DGZ

MACRO PCI33SDGZ
    CLASS PAD ;
    FOREIGN PCI33SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PCI33SDGZ

MACRO PCI66DGZ
    CLASS PAD ;
    FOREIGN PCI66DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PCI66DGZ

MACRO PCI66SDGZ
    CLASS PAD ;
    FOREIGN PCI66SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PCI66SDGZ

MACRO PCORNERDGZ
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN PCORNERDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 246.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE corner ;
    PIN C
        DIRECTION INOUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.000 20.000 150.000 30.000 ;
        RECT  20.000 20.000 30.000 150.000 ;
        RECT  0.000 0.000 150.000 10.000 ;
        RECT  0.000 0.000 10.000 150.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 246.000 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 246.000 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 246.000 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 246.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 246.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 246.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 246.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 246.000 246.000 ;
    END
END PCORNERDGZ

MACRO PDB02DGZ
    CLASS PAD ;
    FOREIGN PDB02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB02DGZ

MACRO PDB02SDGZ
    CLASS PAD ;
    FOREIGN PDB02SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB02SDGZ

MACRO PDB04DGZ
    CLASS PAD ;
    FOREIGN PDB04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB04DGZ

MACRO PDB04SDGZ
    CLASS PAD ;
    FOREIGN PDB04SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB04SDGZ

MACRO PDB08DGZ
    CLASS PAD ;
    FOREIGN PDB08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB08DGZ

MACRO PDB08SDGZ
    CLASS PAD ;
    FOREIGN PDB08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB08SDGZ

MACRO PDB12DGZ
    CLASS PAD ;
    FOREIGN PDB12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB12DGZ

MACRO PDB12SDGZ
    CLASS PAD ;
    FOREIGN PDB12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB12SDGZ

MACRO PDB16DGZ
    CLASS PAD ;
    FOREIGN PDB16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB16DGZ

MACRO PDB16SDGZ
    CLASS PAD ;
    FOREIGN PDB16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB16SDGZ

MACRO PDB24DGZ
    CLASS PAD ;
    FOREIGN PDB24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB24DGZ

MACRO PDB24SDGZ
    CLASS PAD ;
    FOREIGN PDB24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDB24SDGZ

MACRO PDD02DGZ
    CLASS PAD ;
    FOREIGN PDD02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD02DGZ

MACRO PDD02SDGZ
    CLASS PAD ;
    FOREIGN PDD02SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD02SDGZ

MACRO PDD04DGZ
    CLASS PAD ;
    FOREIGN PDD04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD04DGZ

MACRO PDD04SDGZ
    CLASS PAD ;
    FOREIGN PDD04SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD04SDGZ

MACRO PDD08DGZ
    CLASS PAD ;
    FOREIGN PDD08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD08DGZ

MACRO PDD08SDGZ
    CLASS PAD ;
    FOREIGN PDD08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD08SDGZ

MACRO PDD12DGZ
    CLASS PAD ;
    FOREIGN PDD12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD12DGZ

MACRO PDD12SDGZ
    CLASS PAD ;
    FOREIGN PDD12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD12SDGZ

MACRO PDD16DGZ
    CLASS PAD ;
    FOREIGN PDD16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD16DGZ

MACRO PDD16SDGZ
    CLASS PAD ;
    FOREIGN PDD16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD16SDGZ

MACRO PDD24DGZ
    CLASS PAD ;
    FOREIGN PDD24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD24DGZ

MACRO PDD24SDGZ
    CLASS PAD ;
    FOREIGN PDD24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDD24SDGZ

MACRO PDDDGZ
    CLASS PAD ;
    FOREIGN PDDDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  9.395 0.000 35.000 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  0.000 0.000 6.955 246.000 ;
        LAYER VIA12 ;
        RECT  7.400 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA23 ;
        RECT  7.740 245.395 8.610 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA34 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL4 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA45 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL5 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA56 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL6 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA67 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL7 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA78 ;
        RECT  7.635 245.310 8.715 245.670 ;
        LAYER METAL8 ;
        RECT  9.635 0.000 35.000 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  0.000 0.000 6.715 246.000 ;
    END
END PDDDGZ

MACRO PDDSDGZ
    CLASS PAD ;
    FOREIGN PDDSDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  9.395 0.000 35.000 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  0.000 0.000 6.955 246.000 ;
        LAYER VIA12 ;
        RECT  7.400 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA23 ;
        RECT  7.740 245.395 8.610 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA34 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL4 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA45 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL5 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA56 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL6 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA67 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL7 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA78 ;
        RECT  7.635 245.310 8.715 245.670 ;
        LAYER METAL8 ;
        RECT  9.635 0.000 35.000 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  0.000 0.000 6.715 246.000 ;
    END
END PDDSDGZ

MACRO PDDW02DGZ
    CLASS PAD ;
    FOREIGN PDDW02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDDW02DGZ

MACRO PDDW04DGZ
    CLASS PAD ;
    FOREIGN PDDW04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDDW04DGZ

MACRO PDDW08DGZ
    CLASS PAD ;
    FOREIGN PDDW08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDDW08DGZ

MACRO PDDW12DGZ
    CLASS PAD ;
    FOREIGN PDDW12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDDW12DGZ

MACRO PDDW16DGZ
    CLASS PAD ;
    FOREIGN PDDW16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDDW16DGZ

MACRO PDDW24DGZ
    CLASS PAD ;
    FOREIGN PDDW24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDDW24DGZ

MACRO PDDWDGZ
    CLASS PAD ;
    FOREIGN PDDWDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  13.895 0.000 35.000 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  0.000 0.000 6.955 246.000 ;
        LAYER VIA12 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  7.400 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.915 0.740 21.300 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA23 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.915 0.740 21.300 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA34 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL4 ;
        RECT  13.915 0.000 35.000 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA45 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL5 ;
        RECT  13.915 0.000 35.000 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA56 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL6 ;
        RECT  13.915 0.000 35.000 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA67 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL7 ;
        RECT  13.915 0.000 35.000 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA78 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        LAYER METAL8 ;
        RECT  14.135 0.000 35.000 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  0.000 0.000 6.715 246.000 ;
    END
END PDDWDGZ

MACRO PDIDGZ
    CLASS PAD ;
    FOREIGN PDIDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  9.395 0.000 35.000 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  0.000 0.000 6.955 246.000 ;
        LAYER VIA12 ;
        RECT  7.400 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA23 ;
        RECT  7.740 245.395 8.610 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA34 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL4 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA45 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL5 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA56 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL6 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA67 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL7 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA78 ;
        RECT  7.635 245.310 8.715 245.670 ;
        LAYER METAL8 ;
        RECT  9.635 0.000 35.000 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  0.000 0.000 6.715 246.000 ;
    END
END PDIDGZ

MACRO PDISDGZ
    CLASS PAD ;
    FOREIGN PDISDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  9.395 0.000 35.000 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  0.000 0.000 6.955 246.000 ;
        LAYER VIA12 ;
        RECT  7.400 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA23 ;
        RECT  7.740 245.395 8.610 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA34 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL4 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA45 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL5 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA56 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL6 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA67 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL7 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA78 ;
        RECT  7.635 245.310 8.715 245.670 ;
        LAYER METAL8 ;
        RECT  9.635 0.000 35.000 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  0.000 0.000 6.715 246.000 ;
    END
END PDISDGZ

MACRO PDO02CDG
    CLASS PAD ;
    FOREIGN PDO02CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDO02CDG

MACRO PDO04CDG
    CLASS PAD ;
    FOREIGN PDO04CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDO04CDG

MACRO PDO08CDG
    CLASS PAD ;
    FOREIGN PDO08CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDO08CDG

MACRO PDO12CDG
    CLASS PAD ;
    FOREIGN PDO12CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDO12CDG

MACRO PDO16CDG
    CLASS PAD ;
    FOREIGN PDO16CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDO16CDG

MACRO PDO24CDG
    CLASS PAD ;
    FOREIGN PDO24CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDO24CDG

MACRO PDT02DGZ
    CLASS PAD ;
    FOREIGN PDT02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDT02DGZ

MACRO PDT04DGZ
    CLASS PAD ;
    FOREIGN PDT04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDT04DGZ

MACRO PDT08DGZ
    CLASS PAD ;
    FOREIGN PDT08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDT08DGZ

MACRO PDT12DGZ
    CLASS PAD ;
    FOREIGN PDT12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDT12DGZ

MACRO PDT16DGZ
    CLASS PAD ;
    FOREIGN PDT16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDT16DGZ

MACRO PDT24DGZ
    CLASS PAD ;
    FOREIGN PDT24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDT24DGZ

MACRO PDU02DGZ
    CLASS PAD ;
    FOREIGN PDU02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU02DGZ

MACRO PDU02SDGZ
    CLASS PAD ;
    FOREIGN PDU02SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU02SDGZ

MACRO PDU04DGZ
    CLASS PAD ;
    FOREIGN PDU04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU04DGZ

MACRO PDU04SDGZ
    CLASS PAD ;
    FOREIGN PDU04SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU04SDGZ

MACRO PDU08DGZ
    CLASS PAD ;
    FOREIGN PDU08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU08DGZ

MACRO PDU08SDGZ
    CLASS PAD ;
    FOREIGN PDU08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU08SDGZ

MACRO PDU12DGZ
    CLASS PAD ;
    FOREIGN PDU12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU12DGZ

MACRO PDU12SDGZ
    CLASS PAD ;
    FOREIGN PDU12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU12SDGZ

MACRO PDU16DGZ
    CLASS PAD ;
    FOREIGN PDU16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU16DGZ

MACRO PDU16SDGZ
    CLASS PAD ;
    FOREIGN PDU16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU16SDGZ

MACRO PDU24DGZ
    CLASS PAD ;
    FOREIGN PDU24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU24DGZ

MACRO PDU24SDGZ
    CLASS PAD ;
    FOREIGN PDU24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDU24SDGZ

MACRO PDUDGZ
    CLASS PAD ;
    FOREIGN PDUDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  9.395 0.000 35.000 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  0.000 0.000 6.955 246.000 ;
        LAYER VIA12 ;
        RECT  7.400 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA23 ;
        RECT  7.740 245.395 8.610 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA34 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL4 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA45 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL5 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA56 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL6 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA67 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL7 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA78 ;
        RECT  7.635 245.310 8.715 245.670 ;
        LAYER METAL8 ;
        RECT  9.635 0.000 35.000 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  0.000 0.000 6.715 246.000 ;
    END
END PDUDGZ

MACRO PDUSDGZ
    CLASS PAD ;
    FOREIGN PDUSDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  9.395 0.000 35.000 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  0.000 0.000 6.955 246.000 ;
        LAYER VIA12 ;
        RECT  7.400 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA23 ;
        RECT  7.740 245.395 8.610 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA34 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL4 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA45 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL5 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA56 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL6 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA67 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL7 ;
        RECT  9.415 0.000 35.000 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA78 ;
        RECT  7.635 245.310 8.715 245.670 ;
        LAYER METAL8 ;
        RECT  9.635 0.000 35.000 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  0.000 0.000 6.715 246.000 ;
    END
END PDUSDGZ

MACRO PDUW02DGZ
    CLASS PAD ;
    FOREIGN PDUW02DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDUW02DGZ

MACRO PDUW04DGZ
    CLASS PAD ;
    FOREIGN PDUW04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDUW04DGZ

MACRO PDUW08DGZ
    CLASS PAD ;
    FOREIGN PDUW08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDUW08DGZ

MACRO PDUW12DGZ
    CLASS PAD ;
    FOREIGN PDUW12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDUW12DGZ

MACRO PDUW16DGZ
    CLASS PAD ;
    FOREIGN PDUW16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDUW16DGZ

MACRO PDUW24DGZ
    CLASS PAD ;
    FOREIGN PDUW24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PDUW24DGZ

MACRO PDUWDGZ
    CLASS PAD ;
    FOREIGN PDUWDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  13.895 0.000 35.000 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  0.000 0.000 6.955 246.000 ;
        LAYER VIA12 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  7.400 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.915 0.740 21.300 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA23 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.915 0.740 21.300 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA34 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL4 ;
        RECT  13.915 0.000 35.000 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA45 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL5 ;
        RECT  13.915 0.000 35.000 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA56 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL6 ;
        RECT  13.915 0.000 35.000 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA67 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        LAYER METAL7 ;
        RECT  13.915 0.000 35.000 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  0.000 0.000 6.935 246.000 ;
        LAYER VIA78 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        LAYER METAL8 ;
        RECT  14.135 0.000 35.000 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  0.000 0.000 6.715 246.000 ;
    END
END PDUWDGZ

MACRO PDXO01DG
    CLASS PAD ;
    FOREIGN PDXO01DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  56.440 0.000 63.560 0.500 ;
        LAYER METAL3 ;
        RECT  56.440 0.000 63.560 0.500 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  16.440 0.000 23.560 0.500 ;
        LAYER METAL3 ;
        RECT  16.440 0.000 23.560 0.500 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL2 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL3 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL4 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL5 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL6 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL7 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL8 ;
        RECT  46.190 245.000 48.190 246.000 ;
        END
    END XC
    OBS
        LAYER METAL1 ;
        RECT  48.410 0.000 80.000 246.000 ;
        RECT  45.970 0.000 48.410 244.780 ;
        RECT  0.000 0.000 45.970 246.000 ;
        LAYER VIA12 ;
        RECT  46.415 245.395 47.965 245.585 ;
        LAYER METAL2 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  48.430 0.000 56.200 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  23.800 0.000 45.950 246.000 ;
        RECT  16.200 0.740 23.800 246.000 ;
        RECT  0.000 0.000 16.200 246.000 ;
        LAYER VIA23 ;
        RECT  46.755 245.395 47.625 245.585 ;
        LAYER METAL3 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  48.430 0.000 56.200 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  23.800 0.000 45.950 246.000 ;
        RECT  16.200 0.740 23.800 246.000 ;
        RECT  0.000 0.000 16.200 246.000 ;
        LAYER VIA34 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL4 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA45 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL5 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA56 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL6 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA67 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL7 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA78 ;
        RECT  46.650 245.310 47.730 245.670 ;
        LAYER METAL8 ;
        RECT  48.650 0.000 80.000 246.000 ;
        RECT  45.730 0.000 48.650 244.540 ;
        RECT  0.000 0.000 45.730 246.000 ;
    END
END PDXO01DG

MACRO PDXO02DG
    CLASS PAD ;
    FOREIGN PDXO02DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  56.440 0.000 63.560 0.500 ;
        LAYER METAL3 ;
        RECT  56.440 0.000 63.560 0.500 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL2 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL3 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL4 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL5 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL6 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL7 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL8 ;
        RECT  46.190 245.000 48.190 246.000 ;
        END
    END XC
    OBS
        LAYER METAL1 ;
        RECT  48.410 0.000 80.000 246.000 ;
        RECT  45.970 0.000 48.410 244.780 ;
        RECT  0.000 0.000 45.970 246.000 ;
        LAYER VIA12 ;
        RECT  46.415 245.395 47.965 245.585 ;
        LAYER METAL2 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  48.430 0.000 56.200 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA23 ;
        RECT  46.755 245.395 47.625 245.585 ;
        RECT  15.370 0.055 15.970 0.245 ;
        LAYER METAL3 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  48.430 0.000 56.200 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA34 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL4 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA45 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL5 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA56 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL6 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA67 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL7 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA78 ;
        RECT  46.650 245.310 47.730 245.670 ;
        LAYER METAL8 ;
        RECT  48.650 0.000 80.000 246.000 ;
        RECT  45.730 0.000 48.650 244.540 ;
        RECT  0.000 0.000 45.730 246.000 ;
    END
END PDXO02DG

MACRO PDXO03DG
    CLASS PAD ;
    FOREIGN PDXO03DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  56.440 0.000 63.560 0.500 ;
        LAYER METAL3 ;
        RECT  56.440 0.000 63.560 0.500 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL2 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL3 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL4 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL5 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL6 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL7 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL8 ;
        RECT  46.190 245.000 48.190 246.000 ;
        END
    END XC
    OBS
        LAYER METAL1 ;
        RECT  48.410 0.000 80.000 246.000 ;
        RECT  45.970 0.000 48.410 244.780 ;
        RECT  0.000 0.000 45.970 246.000 ;
        LAYER VIA12 ;
        RECT  46.415 245.395 47.965 245.585 ;
        LAYER METAL2 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  48.430 0.000 56.200 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA23 ;
        RECT  46.755 245.395 47.625 245.585 ;
        RECT  15.370 0.055 15.970 0.245 ;
        LAYER METAL3 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  48.430 0.000 56.200 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA34 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL4 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA45 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL5 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA56 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL6 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA67 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL7 ;
        RECT  48.430 0.000 80.000 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA78 ;
        RECT  46.650 245.310 47.730 245.670 ;
        LAYER METAL8 ;
        RECT  48.650 0.000 80.000 246.000 ;
        RECT  45.730 0.000 48.650 244.540 ;
        RECT  0.000 0.000 45.730 246.000 ;
    END
END PDXO03DG

MACRO PDXOE1DG
    CLASS PAD ;
    FOREIGN PDXOE1DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  56.440 0.000 63.560 0.500 ;
        LAYER METAL3 ;
        RECT  56.440 0.000 63.560 0.500 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL2 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL3 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL4 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL5 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL6 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL7 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL8 ;
        RECT  46.190 245.000 48.190 246.000 ;
        END
    END XC
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL2 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL3 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL4 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL5 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL6 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL7 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL8 ;
        RECT  53.390 245.000 55.390 246.000 ;
        END
    END E
    OBS
        LAYER METAL1 ;
        RECT  55.610 0.000 80.000 246.000 ;
        RECT  53.170 0.000 55.610 244.780 ;
        RECT  48.410 0.000 53.170 246.000 ;
        RECT  45.970 0.000 48.410 244.780 ;
        RECT  0.000 0.000 45.970 246.000 ;
        LAYER VIA12 ;
        RECT  53.615 245.395 55.165 245.585 ;
        RECT  46.415 245.395 47.965 245.585 ;
        LAYER METAL2 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  55.630 0.000 56.200 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA23 ;
        RECT  53.955 245.395 54.825 245.585 ;
        RECT  46.755 245.395 47.625 245.585 ;
        RECT  15.370 0.055 15.970 0.245 ;
        LAYER METAL3 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  55.630 0.000 56.200 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA34 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL4 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA45 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL5 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA56 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL6 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA67 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL7 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA78 ;
        RECT  53.850 245.310 54.930 245.670 ;
        RECT  46.650 245.310 47.730 245.670 ;
        LAYER METAL8 ;
        RECT  55.850 0.000 80.000 246.000 ;
        RECT  52.930 0.000 55.850 244.540 ;
        RECT  48.650 0.000 52.930 246.000 ;
        RECT  45.730 0.000 48.650 244.540 ;
        RECT  0.000 0.000 45.730 246.000 ;
    END
END PDXOE1DG

MACRO PDXOE2DG
    CLASS PAD ;
    FOREIGN PDXOE2DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  56.440 0.000 63.560 0.500 ;
        LAYER METAL3 ;
        RECT  56.440 0.000 63.560 0.500 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL2 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL3 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL4 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL5 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL6 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL7 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL8 ;
        RECT  46.190 245.000 48.190 246.000 ;
        END
    END XC
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL2 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL3 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL4 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL5 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL6 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL7 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL8 ;
        RECT  53.390 245.000 55.390 246.000 ;
        END
    END E
    OBS
        LAYER METAL1 ;
        RECT  55.610 0.000 80.000 246.000 ;
        RECT  53.170 0.000 55.610 244.780 ;
        RECT  48.410 0.000 53.170 246.000 ;
        RECT  45.970 0.000 48.410 244.780 ;
        RECT  0.000 0.000 45.970 246.000 ;
        LAYER VIA12 ;
        RECT  53.615 245.395 55.165 245.585 ;
        RECT  46.415 245.395 47.965 245.585 ;
        LAYER METAL2 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  55.630 0.000 56.200 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA23 ;
        RECT  53.955 245.395 54.825 245.585 ;
        RECT  46.755 245.395 47.625 245.585 ;
        RECT  15.370 0.055 15.970 0.245 ;
        LAYER METAL3 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  55.630 0.000 56.200 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA34 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL4 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA45 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL5 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA56 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL6 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA67 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL7 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA78 ;
        RECT  53.850 245.310 54.930 245.670 ;
        RECT  46.650 245.310 47.730 245.670 ;
        LAYER METAL8 ;
        RECT  55.850 0.000 80.000 246.000 ;
        RECT  52.930 0.000 55.850 244.540 ;
        RECT  48.650 0.000 52.930 246.000 ;
        RECT  45.730 0.000 48.650 244.540 ;
        RECT  0.000 0.000 45.730 246.000 ;
    END
END PDXOE2DG

MACRO PDXOE3DG
    CLASS PAD ;
    FOREIGN PDXOE3DG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  56.440 0.000 63.560 0.500 ;
        LAYER METAL3 ;
        RECT  56.440 0.000 63.560 0.500 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL2 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL3 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL4 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL5 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL6 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL7 ;
        RECT  46.190 245.000 48.190 246.000 ;
        LAYER METAL8 ;
        RECT  46.190 245.000 48.190 246.000 ;
        END
    END XC
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL2 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL3 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL4 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL5 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL6 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL7 ;
        RECT  53.390 245.000 55.390 246.000 ;
        LAYER METAL8 ;
        RECT  53.390 245.000 55.390 246.000 ;
        END
    END E
    OBS
        LAYER METAL1 ;
        RECT  55.610 0.000 80.000 246.000 ;
        RECT  53.170 0.000 55.610 244.780 ;
        RECT  48.410 0.000 53.170 246.000 ;
        RECT  45.970 0.000 48.410 244.780 ;
        RECT  0.000 0.000 45.970 246.000 ;
        LAYER VIA12 ;
        RECT  53.615 245.395 55.165 245.585 ;
        RECT  46.415 245.395 47.965 245.585 ;
        LAYER METAL2 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  55.630 0.000 56.200 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA23 ;
        RECT  53.955 245.395 54.825 245.585 ;
        RECT  46.755 245.395 47.625 245.585 ;
        RECT  15.370 0.055 15.970 0.245 ;
        LAYER METAL3 ;
        RECT  63.800 0.000 80.000 246.000 ;
        RECT  56.200 0.740 63.800 246.000 ;
        RECT  55.630 0.000 56.200 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  21.300 0.000 45.950 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  0.000 0.000 13.700 246.000 ;
        LAYER VIA34 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL4 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA45 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL5 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA56 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL6 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA67 ;
        RECT  53.935 245.395 54.845 245.585 ;
        RECT  46.735 245.395 47.645 245.585 ;
        LAYER METAL7 ;
        RECT  55.630 0.000 80.000 246.000 ;
        RECT  53.150 0.000 55.630 244.760 ;
        RECT  48.430 0.000 53.150 246.000 ;
        RECT  45.950 0.000 48.430 244.760 ;
        RECT  0.000 0.000 45.950 246.000 ;
        LAYER VIA78 ;
        RECT  53.850 245.310 54.930 245.670 ;
        RECT  46.650 245.310 47.730 245.670 ;
        LAYER METAL8 ;
        RECT  55.850 0.000 80.000 246.000 ;
        RECT  52.930 0.000 55.850 244.540 ;
        RECT  48.650 0.000 52.930 246.000 ;
        RECT  45.730 0.000 48.650 244.540 ;
        RECT  0.000 0.000 45.730 246.000 ;
    END
END PDXOE3DG

MACRO PFEED0_005Z
    CLASS PAD ;
    FOREIGN PFEED0_005Z 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.005 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 0.005 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 0.005 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 0.005 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 0.005 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 0.005 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 0.005 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 0.005 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 0.005 246.000 ;
    END
END PFEED0_005Z

MACRO PFEED0_01Z
    CLASS PAD ;
    FOREIGN PFEED0_01Z 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.010 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 0.010 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 0.010 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 0.010 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 0.010 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 0.010 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 0.010 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 0.010 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 0.010 246.000 ;
    END
END PFEED0_01Z

MACRO PFEED0_1Z
    CLASS PAD ;
    FOREIGN PFEED0_1Z 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.100 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 0.100 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 0.100 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 0.100 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 0.100 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 0.100 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 0.100 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 0.100 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 0.100 246.000 ;
    END
END PFEED0_1Z

MACRO PFEED10Z
    CLASS PAD ;
    FOREIGN PFEED10Z 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 10.000 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 10.000 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 10.000 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 10.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 10.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 10.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 10.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 10.000 246.000 ;
    END
END PFEED10Z

MACRO PFEED1Z
    CLASS PAD ;
    FOREIGN PFEED1Z 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 1.000 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 1.000 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 1.000 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 1.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 1.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 1.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 1.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 1.000 246.000 ;
    END
END PFEED1Z

MACRO PFEED20Z
    CLASS PAD ;
    FOREIGN PFEED20Z 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 20.000 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 20.000 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 20.000 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 20.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 20.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 20.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 20.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 20.000 246.000 ;
    END
END PFEED20Z

MACRO PFEED5Z
    CLASS PAD ;
    FOREIGN PFEED5Z 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 5.000 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 5.000 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 5.000 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 5.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 5.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 5.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 5.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 5.000 246.000 ;
    END
END PFEED5Z

MACRO PRB08DGZ
    CLASS PAD ;
    FOREIGN PRB08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRB08DGZ

MACRO PRB08SDGZ
    CLASS PAD ;
    FOREIGN PRB08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRB08SDGZ

MACRO PRB12DGZ
    CLASS PAD ;
    FOREIGN PRB12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRB12DGZ

MACRO PRB12SDGZ
    CLASS PAD ;
    FOREIGN PRB12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRB12SDGZ

MACRO PRB16DGZ
    CLASS PAD ;
    FOREIGN PRB16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRB16DGZ

MACRO PRB16SDGZ
    CLASS PAD ;
    FOREIGN PRB16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRB16SDGZ

MACRO PRB24DGZ
    CLASS PAD ;
    FOREIGN PRB24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRB24DGZ

MACRO PRB24SDGZ
    CLASS PAD ;
    FOREIGN PRB24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRB24SDGZ

MACRO PRD08DGZ
    CLASS PAD ;
    FOREIGN PRD08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRD08DGZ

MACRO PRD08SDGZ
    CLASS PAD ;
    FOREIGN PRD08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRD08SDGZ

MACRO PRD12DGZ
    CLASS PAD ;
    FOREIGN PRD12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRD12DGZ

MACRO PRD12SDGZ
    CLASS PAD ;
    FOREIGN PRD12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRD12SDGZ

MACRO PRD16DGZ
    CLASS PAD ;
    FOREIGN PRD16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRD16DGZ

MACRO PRD16SDGZ
    CLASS PAD ;
    FOREIGN PRD16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRD16SDGZ

MACRO PRD24DGZ
    CLASS PAD ;
    FOREIGN PRD24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRD24DGZ

MACRO PRD24SDGZ
    CLASS PAD ;
    FOREIGN PRD24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRD24SDGZ

MACRO PRDW08DGZ
    CLASS PAD ;
    FOREIGN PRDW08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRDW08DGZ

MACRO PRDW12DGZ
    CLASS PAD ;
    FOREIGN PRDW12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRDW12DGZ

MACRO PRDW16DGZ
    CLASS PAD ;
    FOREIGN PRDW16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRDW16DGZ

MACRO PRDW24DGZ
    CLASS PAD ;
    FOREIGN PRDW24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRDW24DGZ

MACRO PRO08CDG
    CLASS PAD ;
    FOREIGN PRO08CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRO08CDG

MACRO PRO12CDG
    CLASS PAD ;
    FOREIGN PRO12CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRO12CDG

MACRO PRO16CDG
    CLASS PAD ;
    FOREIGN PRO16CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRO16CDG

MACRO PRO24CDG
    CLASS PAD ;
    FOREIGN PRO24CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  5.910 0.000 35.000 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  13.700 0.740 21.300 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  5.930 0.000 35.000 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  6.150 0.000 35.000 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRO24CDG

MACRO PRT08DGZ
    CLASS PAD ;
    FOREIGN PRT08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRT08DGZ

MACRO PRT12DGZ
    CLASS PAD ;
    FOREIGN PRT12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRT12DGZ

MACRO PRT16DGZ
    CLASS PAD ;
    FOREIGN PRT16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRT16DGZ

MACRO PRT24DGZ
    CLASS PAD ;
    FOREIGN PRT24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  5.910 0.000 17.075 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 5.465 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  5.930 0.000 13.700 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  5.930 0.000 17.055 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  6.150 0.000 16.835 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRT24DGZ

MACRO PRU08DGZ
    CLASS PAD ;
    FOREIGN PRU08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRU08DGZ

MACRO PRU08SDGZ
    CLASS PAD ;
    FOREIGN PRU08SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRU08SDGZ

MACRO PRU12DGZ
    CLASS PAD ;
    FOREIGN PRU12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRU12DGZ

MACRO PRU12SDGZ
    CLASS PAD ;
    FOREIGN PRU12SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRU12SDGZ

MACRO PRU16DGZ
    CLASS PAD ;
    FOREIGN PRU16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRU16DGZ

MACRO PRU16SDGZ
    CLASS PAD ;
    FOREIGN PRU16SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRU16SDGZ

MACRO PRU24DGZ
    CLASS PAD ;
    FOREIGN PRU24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRU24DGZ

MACRO PRU24SDGZ
    CLASS PAD ;
    FOREIGN PRU24SDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  9.395 0.000 17.075 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.700 0.740 17.055 246.000 ;
        RECT  9.415 0.000 13.700 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  9.415 0.000 17.055 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  9.635 0.000 16.835 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRU24SDGZ

MACRO PRUW08DGZ
    CLASS PAD ;
    FOREIGN PRUW08DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRUW08DGZ

MACRO PRUW12DGZ
    CLASS PAD ;
    FOREIGN PRUW12DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRUW12DGZ

MACRO PRUW16DGZ
    CLASS PAD ;
    FOREIGN PRUW16DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRUW16DGZ

MACRO PRUW24DGZ
    CLASS PAD ;
    FOREIGN PRUW24DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL2 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL3 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL4 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL5 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL6 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL7 ;
        RECT  11.675 245.000 13.675 246.000 ;
        LAYER METAL8 ;
        RECT  11.675 245.000 13.675 246.000 ;
        END
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER METAL2 ;
        RECT  13.940 0.000 21.060 0.500 ;
        LAYER METAL3 ;
        RECT  13.940 0.000 21.060 0.500 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL2 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL3 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL4 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL5 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL6 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL7 ;
        RECT  17.295 245.000 19.295 246.000 ;
        LAYER METAL8 ;
        RECT  17.295 245.000 19.295 246.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL2 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL3 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL4 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL5 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL6 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL7 ;
        RECT  3.690 245.000 5.690 246.000 ;
        LAYER METAL8 ;
        RECT  3.690 245.000 5.690 246.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL2 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL3 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL4 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL5 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL6 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL7 ;
        RECT  7.175 245.000 9.175 246.000 ;
        LAYER METAL8 ;
        RECT  7.175 245.000 9.175 246.000 ;
        END
    END C
    OBS
        LAYER METAL1 ;
        RECT  19.515 0.000 35.000 246.000 ;
        RECT  17.075 0.000 19.515 244.780 ;
        RECT  13.895 0.000 17.075 246.000 ;
        RECT  11.455 0.000 13.895 244.780 ;
        RECT  9.395 0.000 11.455 246.000 ;
        RECT  6.955 0.000 9.395 244.780 ;
        RECT  5.910 0.000 6.955 246.000 ;
        RECT  3.470 0.000 5.910 244.780 ;
        RECT  0.000 0.000 3.470 246.000 ;
        LAYER VIA12 ;
        RECT  17.520 245.395 19.070 245.585 ;
        RECT  11.900 245.395 13.450 245.585 ;
        RECT  3.915 245.395 8.950 245.585 ;
        LAYER METAL2 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA23 ;
        RECT  17.860 245.395 18.730 245.585 ;
        RECT  12.240 245.395 13.110 245.585 ;
        RECT  7.740 245.395 8.610 245.585 ;
        RECT  4.255 245.395 5.125 245.585 ;
        LAYER METAL3 ;
        RECT  21.300 0.000 35.000 246.000 ;
        RECT  19.535 0.740 21.300 246.000 ;
        RECT  17.055 0.740 19.535 244.760 ;
        RECT  13.915 0.740 17.055 246.000 ;
        RECT  13.700 0.740 13.915 244.760 ;
        RECT  11.435 0.000 13.700 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA34 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL4 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA45 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL5 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA56 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL6 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA67 ;
        RECT  17.840 245.395 18.750 245.585 ;
        RECT  12.220 245.395 13.130 245.585 ;
        RECT  7.720 245.395 8.630 245.585 ;
        RECT  4.235 245.395 5.145 245.585 ;
        LAYER METAL7 ;
        RECT  19.535 0.000 35.000 246.000 ;
        RECT  17.055 0.000 19.535 244.760 ;
        RECT  13.915 0.000 17.055 246.000 ;
        RECT  11.435 0.000 13.915 244.760 ;
        RECT  9.415 0.000 11.435 246.000 ;
        RECT  6.935 0.000 9.415 244.760 ;
        RECT  5.930 0.000 6.935 246.000 ;
        RECT  3.450 0.000 5.930 244.760 ;
        RECT  0.000 0.000 3.450 246.000 ;
        LAYER VIA78 ;
        RECT  17.755 245.310 18.835 245.670 ;
        RECT  12.135 245.310 13.215 245.670 ;
        RECT  7.635 245.310 8.715 245.670 ;
        RECT  4.150 245.310 5.230 245.670 ;
        LAYER METAL8 ;
        RECT  19.755 0.000 35.000 246.000 ;
        RECT  16.835 0.000 19.755 244.540 ;
        RECT  14.135 0.000 16.835 246.000 ;
        RECT  11.215 0.000 14.135 244.540 ;
        RECT  9.635 0.000 11.215 246.000 ;
        RECT  6.715 0.000 9.635 244.540 ;
        RECT  6.150 0.000 6.715 246.000 ;
        RECT  3.230 0.000 6.150 244.540 ;
        RECT  0.000 0.000 3.230 246.000 ;
    END
END PRUW24DGZ

MACRO PVDD1DGZ
    CLASS PAD POWER ;
    FOREIGN PVDD1DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        CLASS CORE ;
        LAYER METAL2 ;
        RECT  4.180 241.940 30.820 246.000 ;
        LAYER METAL3 ;
        RECT  4.180 241.940 30.820 246.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL2 ;
        RECT  31.420 0.000 35.000 246.000 ;
        RECT  3.580 0.000 31.420 241.340 ;
        RECT  0.000 0.000 3.580 246.000 ;
        LAYER VIA23 ;
        RECT  4.380 241.945 30.490 243.755 ;
        LAYER METAL3 ;
        RECT  31.420 0.000 35.000 246.000 ;
        RECT  3.580 0.000 31.420 241.340 ;
        RECT  0.000 0.000 3.580 246.000 ;
        LAYER VIA34 ;
        RECT  4.435 242.420 29.825 243.510 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 35.000 246.000 ;
    END
END PVDD1DGZ

MACRO PVDD2DGZ
    CLASS PAD ;
    FOREIGN PVDD2DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 35.000 246.000 ;
    END
END PVDD2DGZ

MACRO PVDD2POC
    CLASS PAD ;
    FOREIGN PVDD2POC 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 35.000 246.000 ;
    END
END PVDD2POC

MACRO PVSS1DGZ
    CLASS PAD POWER ;
    FOREIGN PVSS1DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        CLASS CORE ;
        LAYER METAL2 ;
        RECT  4.180 239.190 30.820 246.000 ;
        LAYER METAL3 ;
        RECT  4.180 239.190 30.820 246.000 ;
        END
    END VSS
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL2 ;
        RECT  31.420 0.000 35.000 246.000 ;
        RECT  3.580 0.000 31.420 238.590 ;
        RECT  0.000 0.000 3.580 246.000 ;
        LAYER METAL3 ;
        RECT  31.420 0.000 35.000 246.000 ;
        RECT  3.580 0.000 31.420 238.590 ;
        RECT  0.000 0.000 3.580 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 35.000 246.000 ;
    END
END PVSS1DGZ

MACRO PVSS2DGZ
    CLASS PAD ;
    FOREIGN PVSS2DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL2 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL3 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 35.000 246.000 ;
    END
END PVSS2DGZ

MACRO PVSS3DGZ
    CLASS PAD ;
    FOREIGN PVSS3DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 246.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        CLASS CORE ;
        LAYER METAL2 ;
        RECT  5.280 238.140 29.720 246.000 ;
        LAYER METAL3 ;
        RECT  5.280 238.140 29.720 246.000 ;
        END
    END VSS
    OBS
        LAYER METAL1 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL2 ;
        RECT  30.320 0.000 35.000 246.000 ;
        RECT  4.680 0.000 30.320 237.540 ;
        RECT  0.000 0.000 4.680 246.000 ;
        LAYER METAL3 ;
        RECT  30.320 0.000 35.000 246.000 ;
        RECT  4.680 0.000 30.320 237.540 ;
        RECT  0.000 0.000 4.680 246.000 ;
        LAYER METAL4 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL5 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL6 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL7 ;
        RECT  0.000 0.000 35.000 246.000 ;
        LAYER METAL8 ;
        RECT  0.000 0.000 35.000 246.000 ;
    END
END PVSS3DGZ

END LIBRARY
