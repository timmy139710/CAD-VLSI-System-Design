#******
# Preview export LEF
#
#        Preview sub-version 4.4.2.100.41
#
# TECH LIB NAME: tsmc13
#
# RC values have been extracted from TSMC's worst case interconnect
# tables included with CL013G FSG spice model version 1.3P1.
# Document No. T-013-LO-SP-004-PR Rev1.3P1 Jan. 15, 2002
# RC values are also compatible with CL013LV FSG version 1.1
# Document No. T-013-LO-SP-009 Rev1.1 Jan. 29, 2002
#
# Resistance and Capacitance Values
# ---------------------------------
# The LEF technology files included in this directory contain resistance and
# capacitance (RC) values for the purpose of timing driven place & route.
# Please note that the RC values contained in this tech file were created using
# the worst case interconnect models from the foundry and assume a full metal
# route at every grid location on every metal layer, so the values are
# intentionally very conservative. It is assumed that this technology file will
# be used only as a starting point for creating initial timing driven place &
# route runs during the development of your own more accurate RC values,
# tailored to your specific place & route environment. AS A RESULT, TIMING
# NUMBERS DERIVED FROM THESE RC VALUES MAY BE SIGNIFICANTLY SLOWER THAN
# REALITY.
# 
# The RC values used in the LEF technology file are to be used only for timing
# driven place & route. Due to accuracy limitations, please do not attempt to
# use this file for chip-level RC extraction in conjunction with your sign-off
# timing simulations. For chip-level extraction, please use a dedicated
# extraction tool such as HyperExtract, starRC or Simplex, etc.
#
# Antenna Effect Properties
# -------------------------
# Antenna effect properties were modeled based on the following design rule
# document:
#
# Document No. T-013-LO-DR-001 (TSMC 0.13um Logic 1P8M Salicide 1.0V/2.5V,
#                            1.2V/2.5V, 1.0V/3.3V, 1.2V/3.3V Design Rule
#                            version 1.5 8/1/02 )
#
# DO NOT USE SILICON ENSEMBLE OR WROUTE AS A SIGN-OFF VALIDATION FLOW FOR
# PROCESS ANTENNA EFFECT VIOLATIONS.  Foundry DRC command files should always be
# used for sign-off validation of process antenna effect in your design.
#
# $Id: tsmc13fsg_8lm_tech.lef,v 1.3 2004-03-05 19:15:54-08 wching Exp $
#
#******

##############################
# Modified by CIC 2005/07/29 #
##############################
VERSION 5.5 ;
##############################
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;

UNITS
    DATABASE MICRONS 2000  ;
END UNITS

MANUFACTURINGGRID 0.005 ;
USEMINSPACING OBS OFF ;

LAYER POLY1
    TYPE MASTERSLICE ;
END POLY1

LAYER METAL1
    TYPE ROUTING ;
    WIDTH 0.160 ;
    SPACING 0.180 ;
    SPACING 0.18 LENGTHTHRESHOLD  1.0 ;
    SPACING 0.22 RANGE 0.3 10.0 USELENGTHTHRESHOLD ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.410 ;
    OFFSET 0.205 ;
    DIRECTION HORIZONTAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.122 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.26 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL1 = 0.117 ohm/sq) = 1.1700e-01
    RESISTANCE RPERSQ      1.1700e-01 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M2-M1-PO1(FOX):0.16:0.18: CAP1 = (Cb_a * PO1(FOX) ratio + Ct_a * M2 ratio) / M1 width = 0.0761773073136342
      # M2-M1-PO1(FOX):0.16:0.18: CAP1 = (6.44e-03 * 1 + 1.11e-02 * 0.401752173913043) / 0.14308 = 0.0761773073136342
      # M3-M1-PO1(FOX):0.16:0.18: CAP2 = (Cb_a * PO1(FOX) ratio + Ct_a * M3 ratio) / M1 width = 0.0163485392787252
      # M3-M1-PO1(FOX):0.16:0.18: CAP2 = (6.44e-03 * 0 + 3.91e-03 * 0.598247826086957) / 0.14308 = 0.0163485392787252
      # CAP = (0.0761773073136342 + 0.0163485392787252) * 0.001 pF/fF = 9.2526e-05
    CAPACITANCE CPERSQDIST 9.2526e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M2-M1-PO1(FOX):0.16:0.18: ECAP1 = Cfb * PO1(FOX) ratio + Cft * M2 ratio = 0.019456896
      # M2-M1-PO1(FOX):0.16:0.18: ECAP1 = 1.65e-02 * 1 + 7.36e-03 * 0.401752173913043 = 0.019456896
      # M3-M1-PO1(FOX):0.16:0.18: ECAP2 = Cfb * PO1(FOX) ratio + Cft * M3 ratio = 0.00176483108695652
      # M3-M1-PO1(FOX):0.16:0.18: ECAP2 = 1.71e-02 * 0 + 2.95e-03 * 0.598247826086957 = 0.00176483108695652
      # M3-M1-PO1(FOX):0.16:0.18: Cc = 7.88e-02
      # ECAP = (0.019456896 + 0.00176483108695652 + 7.88e-02) * 0.001 pF/fF = 1.0002e-04
    EDGECAPACITANCE        1.0002e-04 ;
END METAL1

LAYER VIA12
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA12

LAYER METAL2
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.460 ;
    OFFSET 0.230 ;
    DIRECTION VERTICAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL2 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M3-M2-M1:0.2:0.21: CAP1 = (Cb_a * M1 ratio + Ct_a * M3 ratio) / M2 width = 0.073567268827456
      # M3-M2-M1:0.2:0.21: CAP1 = (1.43e-02 * 0.5 + 1.43e-02 * 0.450746341463415) / 0.184806 = 0.073567268827456
      # M4-M2-PO1(FOX):0.2:0.21: CAP2 = (Cb_a * PO1(FOX) ratio + Ct_a * M4 ratio) / M2 width = 0.03232433457577
      # M4-M2-PO1(FOX):0.2:0.21: CAP2 = (6.40e-03 * 0.5 + 5.05e-03 * 0.549253658536585) / 0.184806 = 0.03232433457577
      # CAP = (0.073567268827456 + 0.03232433457577) * 0.001 pF/fF = 1.0589e-04
    CAPACITANCE CPERSQDIST 1.0589e-04 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M3-M2-M1:0.2:0.21: ECAP1 = Cfb * M1 ratio + Cft * M3 ratio = 0.00782774687804878
      # M3-M2-M1:0.2:0.21: ECAP1 = 8.11e-03 * 0.5 + 8.37e-03 * 0.450746341463415 = 0.00782774687804878
      # M4-M2-PO1(FOX):0.2:0.21: ECAP2 = Cfb * PO1(FOX) ratio + Cft * M4 ratio = 0.00411886541463415
      # M4-M2-PO1(FOX):0.2:0.21: ECAP2 = 4.36e-03 * 0.5 + 3.53e-03 * 0.549253658536585 = 0.00411886541463415
      # M4-M2-PO1(FOX):0.2:0.21: Cc = 8.65e-02
      # ECAP = (0.00782774687804878 + 0.00411886541463415 + 8.65e-02) * 0.001 pF/fF = 9.8447e-05
    EDGECAPACITANCE        9.8447e-05 ;
END METAL2

LAYER VIA23
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA23

LAYER METAL3
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.410 ;
    OFFSET 0.205 ;
    DIRECTION HORIZONTAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL3 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M4-M3-M2:0.2:0.21: CAP1 = (Cb_a * M2 ratio + Ct_a * M4 ratio) / M3 width = 0.0621739130434783
      # M4-M3-M2:0.2:0.21: CAP1 = (1.43e-02 * 0.401752173913043 + 1.43e-02 * 0.401752173913043) / 0.184806 = 0.0621739130434783
      # M5-M3-M1:0.2:0.21: CAP2 = (Cb_a * M1 ratio + Ct_a * M5 ratio) / M3 width = 0.0326953835020414
      # M5-M3-M1:0.2:0.21: CAP2 = (5.05e-03 * 0.598247826086957 + 5.05e-03 * 0.598247826086957) / 0.184806 = 0.0326953835020414
      # CAP = (0.0621739130434783 + 0.0326953835020414) * 0.001 pF/fF = 9.4869e-05
    CAPACITANCE CPERSQDIST 9.4869e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M4-M3-M2:0.2:0.21: ECAP1 = Cfb * M2 ratio + Cft * M4 ratio = 0.00662087582608696
      # M4-M3-M2:0.2:0.21: ECAP1 = 8.11e-03 * 0.401752173913043 + 8.37e-03 * 0.401752173913043 = 0.00662087582608696
      # M5-M3-M1:0.2:0.21: ECAP2 = Cfb * M1 ratio + Cft * M5 ratio = 0.00433729673913043
      # M5-M3-M1:0.2:0.21: ECAP2 = 3.63e-03 * 0.598247826086957 + 3.62e-03 * 0.598247826086957 = 0.00433729673913043
      # M5-M3-M1:0.2:0.21: Cc = 8.70e-02
      # ECAP = (0.00662087582608696 + 0.00433729673913043 + 8.70e-02) * 0.001 pF/fF = 9.7958e-05
    EDGECAPACITANCE        9.7958e-05 ;
END METAL3

LAYER VIA34
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA34

LAYER METAL4
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.460 ;
    OFFSET 0.230 ;
    DIRECTION VERTICAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL4 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M5-M4-M3:0.2:0.21: CAP1 = (Cb_a * M3 ratio + Ct_a * M5 ratio) / M4 width = 0.0697560975609756
      # M5-M4-M3:0.2:0.21: CAP1 = (1.43e-02 * 0.450746341463415 + 1.43e-02 * 0.450746341463415) / 0.184806 = 0.0697560975609756
      # M6-M4-M2:0.2:0.21: CAP2 = (Cb_a * M2 ratio + Ct_a * M6 ratio) / M4 width = 0.0300177588997084
      # M6-M4-M2:0.2:0.21: CAP2 = (5.05e-03 * 0.549253658536585 + 5.05e-03 * 0.549253658536585) / 0.184806 = 0.0300177588997084
      # CAP = (0.0697560975609756 + 0.0300177588997084) * 0.001 pF/fF = 9.9774e-05
    CAPACITANCE CPERSQDIST 9.9774e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M5-M4-M3:0.2:0.21: ECAP1 = Cfb * M3 ratio + Cft * M5 ratio = 0.00742829970731707
      # M5-M4-M3:0.2:0.21: ECAP1 = 8.11e-03 * 0.450746341463415 + 8.37e-03 * 0.450746341463415 = 0.00742829970731707
      # M6-M4-M2:0.2:0.21: ECAP2 = Cfb * M2 ratio + Cft * M6 ratio = 0.00398208902439024
      # M6-M4-M2:0.2:0.21: ECAP2 = 3.63e-03 * 0.549253658536585 + 3.62e-03 * 0.549253658536585 = 0.00398208902439024
      # M6-M4-M2:0.2:0.21: Cc = 8.70e-02
      # ECAP = (0.00742829970731707 + 0.00398208902439024 + 8.70e-02) * 0.001 pF/fF = 9.8410e-05
    EDGECAPACITANCE        9.8410e-05 ;
END METAL4

LAYER VIA45
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA45

LAYER METAL5
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.410 ;
    OFFSET 0.205 ;
    DIRECTION HORIZONTAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL5 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M6-M5-M4:0.2:0.21: CAP1 = (Cb_a * M4 ratio + Ct_a * M6 ratio) / M5 width = 0.0621739130434783
      # M6-M5-M4:0.2:0.21: CAP1 = (1.43e-02 * 0.401752173913043 + 1.43e-02 * 0.401752173913043) / 0.184806 = 0.0621739130434783
      # M7-M5-M3:0.2:0.21: CAP2 = (Cb_a * M3 ratio + Ct_a * M7 ratio) / M5 width = 0.0326953835020414
      # M7-M5-M3:0.2:0.21: CAP2 = (5.05e-03 * 0.598247826086957 + 5.05e-03 * 0.598247826086957) / 0.184806 = 0.0326953835020414
      # CAP = (0.0621739130434783 + 0.0326953835020414) * 0.001 pF/fF = 9.4869e-05
    CAPACITANCE CPERSQDIST 9.4869e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M6-M5-M4:0.2:0.21: ECAP1 = Cfb * M4 ratio + Cft * M6 ratio = 0.00662087582608696
      # M6-M5-M4:0.2:0.21: ECAP1 = 8.11e-03 * 0.401752173913043 + 8.37e-03 * 0.401752173913043 = 0.00662087582608696
      # M7-M5-M3:0.2:0.21: ECAP2 = Cfb * M3 ratio + Cft * M7 ratio = 0.00433729673913043
      # M7-M5-M3:0.2:0.21: ECAP2 = 3.63e-03 * 0.598247826086957 + 3.62e-03 * 0.598247826086957 = 0.00433729673913043
      # M7-M5-M3:0.2:0.21: Cc = 8.70e-02
      # ECAP = (0.00662087582608696 + 0.00433729673913043 + 8.70e-02) * 0.001 pF/fF = 9.7958e-05
    EDGECAPACITANCE        9.7958e-05 ;
END METAL5

LAYER VIA56
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA56

LAYER METAL6
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.460 ;
    OFFSET 0.230 ;
    DIRECTION VERTICAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL6 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M7-M6-M5:0.2:0.21: CAP1 = (Cb_a * M5 ratio + Ct_a * M7 ratio) / M6 width = 0.058130081300813
      # M7-M6-M5:0.2:0.21: CAP1 = (1.43e-02 * 0.450746341463415 + 1.43e-02 * 0.30049756097561) / 0.184806 = 0.058130081300813
      # M8-M6-M4:0.2:0.21: CAP2 = (Cb_a * M4 ratio + Ct_a * M8 ratio) / M6 width = 0.0322687688579428
      # M8-M6-M4:0.2:0.21: CAP2 = (5.05e-03 * 0.549253658536585 + 4.56e-03 * 0.69950243902439) / 0.184806 = 0.0322687688579428
      # CAP = (0.058130081300813 + 0.0322687688579428) * 0.001 pF/fF = 9.0399e-05
    CAPACITANCE CPERSQDIST 9.0399e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M7-M6-M5:0.2:0.21: ECAP1 = Cfb * M5 ratio + Cft * M7 ratio = 0.00617071741463415
      # M7-M6-M5:0.2:0.21: ECAP1 = 8.11e-03 * 0.450746341463415 + 8.37e-03 * 0.30049756097561 = 0.00617071741463415
      # M8-M6-M4:0.2:0.21: ECAP2 = Cfb * M4 ratio + Cft * M8 ratio = 0.00442002941463415
      # M8-M6-M4:0.2:0.21: ECAP2 = 3.73e-03 * 0.549253658536585 + 3.39e-03 * 0.69950243902439 = 0.00442002941463415
      # M8-M6-M4:0.2:0.21: Cc = 8.73e-02
      # ECAP = (0.00617071741463415 + 0.00442002941463415 + 8.73e-02) * 0.001 pF/fF = 9.7891e-05
    EDGECAPACITANCE        9.7891e-05 ;
END METAL6

LAYER VIA67
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA67

LAYER METAL7
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.615 ;
    OFFSET 0.205 ;
    DIRECTION HORIZONTAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL7 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M8-M7-M6:0.2:0.41: CAP1 = (Cb_a * M6 ratio + Ct_a * M8 ratio) / M7 width = 0.0521304244309779
      # M8-M7-M6:0.2:0.41: CAP1 = (1.43e-02 * 0.401752173913043 + 1.10e-02 * 0.353541739130435) / 0.184806 = 0.0521304244309779
      # M7-M5:0.2:0.41: CAP2 = Ca * M5 ratio / M7 width = 0.0163476917510207
      # M7-M5:0.2:0.41: CAP2 = 5.05e-03 * 0.598247826086957 / 0.184806 = 0.0163476917510207
      # CAP = (0.0521304244309779 + 0.0163476917510207) * 0.001 pF/fF = 6.8478e-05
    CAPACITANCE CPERSQDIST 6.8478e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M8-M7-M6:0.2:0.41: ECAP1 = Cfb * M6 ratio + Cft * M8 ratio = 0.00965490626086957
      # M8-M7-M6:0.2:0.41: ECAP1 = 1.40e-02 * 0.401752173913043 + 1.14e-02 * 0.353541739130435 = 0.00965490626086957
      # M7-M5:0.2:0.41: ECAP2 = Cf * M5 ratio = 0.00506715908695652
      # M7-M5:0.2:0.41: ECAP2 = 8.47e-03 * 0.598247826086957 = 0.00506715908695652
      # M7-M5:0.2:0.41: Cc = 5.33e-02
      # ECAP = (0.00965490626086957 + 0.00506715908695652 + 5.33e-02) * 0.001 pF/fF = 6.8022e-05
    EDGECAPACITANCE        6.8022e-05 ;
END METAL7

LAYER VIA78
    TYPE CUT ;
    SPACING 0.350 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA78

LAYER METAL8
    TYPE ROUTING ;
    WIDTH 0.440 ;
    SPACING 0.460 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 1.150 ;
    OFFSET 0.230 ;
    DIRECTION VERTICAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.562 ;
    MINIMUMCUT 2 WIDTH 1.80 ;
    THICKNESS 0.90 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 51270 ) ( 1 57980 ) ) ;
      # (Worst case resistance model for METAL8 = 0.027 ohm/sq) = 2.7000e-02
    RESISTANCE RPERSQ      2.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M8-M7:0.44:0.66: CAP1 = Ca * M7 ratio / M8 width = 0.0178861876602966
      # M8-M7:0.44:0.66: CAP1 = 2.42e-02 * 0.30049756097561 / 0.406573 = 0.0178861876602966
      # M8-M6:0.44:0.66: CAP2 = Ca * M6 ratio / M8 width = 0.0172048424028253
      # M8-M6:0.44:0.66: CAP2 = 1.00e-02 * 0.69950243902439 / 0.406573 = 0.0172048424028253
      # CAP = (0.0178861876602966 + 0.0172048424028253) * 0.001 pF/fF = 3.5091e-05
    CAPACITANCE CPERSQDIST 3.5091e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M8-M7:0.44:0.66: ECAP1 = Cf * M7 ratio = 0.00558925463414634
      # M8-M7:0.44:0.66: ECAP1 = 1.86e-02 * 0.30049756097561 = 0.00558925463414634
      # M8-M6:0.44:0.66: ECAP2 = Cf * M6 ratio = 0.00647739258536585
      # M8-M6:0.44:0.66: ECAP2 = 9.26e-03 * 0.69950243902439 = 0.00647739258536585
      # M8-M6:0.44:0.66: Cc = 7.25e-02
      # ECAP = (0.00558925463414634 + 0.00647739258536585 + 7.25e-02) * 0.001 pF/fF = 8.4567e-05
    EDGECAPACITANCE        8.4567e-05 ;
END METAL8

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIARULE VIA1ARRAY GENERATE
    LAYER METAL1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA1ARRAY

VIARULE VIA2ARRAY GENERATE
    LAYER METAL2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA2ARRAY

VIARULE VIA3ARRAY GENERATE
    LAYER METAL3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA3ARRAY

VIARULE VIA4ARRAY GENERATE
    LAYER METAL4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA4ARRAY

VIARULE VIA5ARRAY GENERATE
    LAYER METAL5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA5ARRAY

VIARULE VIA6ARRAY GENERATE
    LAYER METAL6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL7 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA6ARRAY

VIARULE VIA7ARRAY GENERATE
    LAYER METAL7 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL8 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER VIA78 ;
        RECT -0.180 -0.180 0.180 0.180 ;
        SPACING 0.900 BY 0.900 ;
END VIA7ARRAY

VIARULE TURNM1 GENERATE
    LAYER METAL1 ;
        DIRECTION VERTICAL ;

    LAYER METAL1 ;
        DIRECTION HORIZONTAL ;
END TURNM1

VIARULE TURNM2 GENERATE
    LAYER METAL2 ;
        DIRECTION VERTICAL ;

    LAYER METAL2 ;
        DIRECTION HORIZONTAL ;
END TURNM2

VIARULE TURNM3 GENERATE
    LAYER METAL3 ;
        DIRECTION VERTICAL ;

    LAYER METAL3 ;
        DIRECTION HORIZONTAL ;
END TURNM3

VIARULE TURNM4 GENERATE
    LAYER METAL4 ;
        DIRECTION VERTICAL ;

    LAYER METAL4 ;
        DIRECTION HORIZONTAL ;
END TURNM4

VIARULE TURNM5 GENERATE
    LAYER METAL5 ;
        DIRECTION VERTICAL ;

    LAYER METAL5 ;
        DIRECTION HORIZONTAL ;
END TURNM5

VIARULE TURNM6 GENERATE
    LAYER METAL6 ;
        DIRECTION VERTICAL ;

    LAYER METAL6 ;
        DIRECTION HORIZONTAL ;
END TURNM6

VIARULE TURNM7 GENERATE
    LAYER METAL7 ;
        DIRECTION VERTICAL ;

    LAYER METAL7 ;
        DIRECTION HORIZONTAL ;
END TURNM7

VIARULE TURNM8 GENERATE
    LAYER METAL8 ;
        DIRECTION VERTICAL ;

    LAYER METAL8 ;
        DIRECTION HORIZONTAL ;
END TURNM8

SPACING
    SAMENET METAL1 METAL1 0.180  ;
    SAMENET METAL2 METAL2 0.210  STACK ;
    SAMENET METAL3 METAL3 0.210  STACK ;
    SAMENET METAL4 METAL4 0.210  STACK ;
    SAMENET METAL5 METAL5 0.210  STACK ;
    SAMENET METAL6 METAL6 0.210  STACK ;
    SAMENET METAL7 METAL7 0.210  STACK ;
    SAMENET METAL8 METAL8 0.460  ;
    SAMENET VIA12 VIA12 0.220  ;
    SAMENET VIA23 VIA23 0.220  ;
    SAMENET VIA34 VIA34 0.220  ;
    SAMENET VIA45 VIA45 0.220  ;
    SAMENET VIA56 VIA56 0.220  ;
    SAMENET VIA67 VIA67 0.220  ;
    SAMENET VIA78 VIA78 0.350  ;
    SAMENET VIA12 VIA23 0.0 STACK ;
    SAMENET VIA23 VIA34 0.0 STACK ;
    SAMENET VIA34 VIA45 0.0 STACK ;
    SAMENET VIA45 VIA56 0.0 STACK ;
    SAMENET VIA56 VIA67 0.0 STACK ;
    SAMENET VIA67 VIA78 0.0 STACK ;
END SPACING

VIA VIA12_H DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL1 ;
        RECT -0.145 -0.105 0.145 0.105 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA12_H

VIA VIA12_V DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL1 ;
        RECT -0.105 -0.145 0.105 0.145 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA12_V

VIA VIA12_X DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL1 ;
        RECT -0.145 -0.105 0.145 0.105 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA12_X

VIA VIA12_XR DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL1 ;
        RECT -0.105 -0.145 0.105 0.145 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA12_XR

VIA VIA23_H DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA23_H

VIA VIA23_V DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA23_V

VIA VIA23_X DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA23_X

VIA VIA23_XR DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA23_XR

VIA VIA34_H DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA34_H

VIA VIA34_V DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA34_V

VIA VIA34_X DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA34_X

VIA VIA34_XR DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA34_XR

VIA VIA45_H DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA45_H

VIA VIA45_V DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA45_V

VIA VIA45_X DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA45_X

VIA VIA45_XR DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA45_XR

VIA VIA56_H DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA56_H

VIA VIA56_V DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA56_V

VIA VIA56_X DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA56_X

VIA VIA56_XR DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA56_XR

VIA VIA67_H DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA67_H

VIA VIA67_V DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA67_V

VIA VIA67_X DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA67_X

VIA VIA67_XR DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA67_XR

VIA VIA78_H DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 6.3000e-01
    RESISTANCE 6.3000e-01 ;
    LAYER METAL7 ;
        RECT -0.23 -0.19 0.23 0.19 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 0.27 0.27 ;
END VIA78_H

VIA VIA78_V DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 6.3000e-01
    RESISTANCE 6.3000e-01 ;
    LAYER METAL7 ;
        RECT -0.19 -0.23 0.19 0.23 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 0.27 0.27 ;
END VIA78_V

VIA VIA78_XR DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 6.3000e-01
    RESISTANCE 6.3000e-01 ;
    LAYER METAL7 ;
        RECT -0.19 -0.23 0.19 0.23 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 0.27 0.27 ;
END VIA78_XR

VIA VIA23_TOS DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.1 -0.370 0.1 0.370 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA23_TOS

VIA VIA34_TOS_E DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.580 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA34_TOS_E

VIA VIA34_TOS_W DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.580 -0.1 0.145 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA34_TOS_W

VIA VIA45_TOS DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.1 -0.370 0.1 0.370 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA45_TOS

VIA VIA56_TOS_E DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.580 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA56_TOS_E

VIA VIA56_TOS_W DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.580 -0.1 0.145 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA56_TOS_W

VIA VIA67_TOS DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.1 -0.370 0.1 0.370 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA67_TOS

VIA VIA12_2CUT_E DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL1 ;
        RECT -0.145 -0.105 0.625 0.105 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA12_2CUT_E

VIA VIA12_2CUT_W DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL1 ;
        RECT -0.625 -0.105 0.145 0.105 ;
    LAYER VIA12 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA12_2CUT_W

VIA VIA12_2CUT_N DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL1 ;
        RECT -0.105 -0.145 0.105 0.625 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA12_2CUT_N

VIA VIA12_2CUT_S DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL1 ;
        RECT -0.105 -0.625 0.105 0.145 ;
    LAYER VIA12 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA12_2CUT_S

VIA VIA23_2CUT_E DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA23_2CUT_E

VIA VIA23_2CUT_W DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL2 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA23 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA23_2CUT_W

VIA VIA23_2CUT_N DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA23_2CUT_N

VIA VIA23_2CUT_S DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL2 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA23 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA23_2CUT_S

VIA VIA34_2CUT_E DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA34_2CUT_E

VIA VIA34_2CUT_W DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL3 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA34 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA34_2CUT_W

VIA VIA34_2CUT_N DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA34_2CUT_N

VIA VIA34_2CUT_S DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL3 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA34 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA34_2CUT_S

VIA VIA45_2CUT_E DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA45_2CUT_E

VIA VIA45_2CUT_W DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL4 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA45 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA45_2CUT_W

VIA VIA45_2CUT_N DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA45_2CUT_N

VIA VIA45_2CUT_S DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL4 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA45 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA45_2CUT_S

VIA VIA56_2CUT_E DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA56_2CUT_E

VIA VIA56_2CUT_W DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL5 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA56 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA56_2CUT_W

VIA VIA56_2CUT_N DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA56_2CUT_N

VIA VIA56_2CUT_S DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL5 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA56 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA56_2CUT_S

VIA VIA67_2CUT_E DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL7 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA67_2CUT_E

VIA VIA67_2CUT_W DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL6 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA67 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA67_2CUT_W

VIA VIA67_2CUT_N DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL7 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA67_2CUT_N

VIA VIA67_2CUT_S DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL6 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA67 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA67_2CUT_S

VIA VIA78_2CUT_E DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 3.1500e-01
    RESISTANCE 3.1500e-01 ;
    LAYER METAL7 ;
        RECT -0.23 -0.19 1.13 0.19 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        RECT 0.72 -0.18 1.08 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 1.17 0.27 ;
END VIA78_2CUT_E

VIA VIA78_2CUT_W DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 3.1500e-01
    RESISTANCE 3.1500e-01 ;
    LAYER METAL7 ;
        RECT -1.13 -0.19 0.23 0.19 ;
    LAYER VIA78 ;
        RECT -1.08 -0.18 -0.72 0.18 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -1.17 -0.27 0.27 0.27 ;
END VIA78_2CUT_W

VIA VIA78_2CUT_N DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 3.1500e-01
    RESISTANCE 3.1500e-01 ;
    LAYER METAL7 ;
        RECT -0.19 -0.23 0.19 1.13 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        RECT -0.18 0.72 0.18 1.08 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 0.27 1.17 ;
END VIA78_2CUT_N

VIA VIA78_2CUT_S DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 3.1500e-01
    RESISTANCE 3.1500e-01 ;
    LAYER METAL7 ;
        RECT -0.19 -1.13 0.19 0.23 ;
    LAYER VIA78 ;
        RECT -0.18 -1.08 0.18 -0.72 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -1.17 0.27 0.27 ;
END VIA78_2CUT_S

SITE TSM13SITE
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.460 BY 3.690 ;
END TSM13SITE

MACRO FILL64
    CLASS CORE SPACER ;
    FOREIGN FILL64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 29.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 29.440 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 29.440 3.940 ;
        END
    END VDD
END FILL64

MACRO FILL32
    CLASS CORE SPACER ;
    FOREIGN FILL32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 14.720 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 14.720 3.940 ;
        END
    END VDD
END FILL32

MACRO FILL16
    CLASS CORE SPACER ;
    FOREIGN FILL16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 7.360 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 7.360 3.940 ;
        END
    END VDD
END FILL16

MACRO FILL8
    CLASS CORE SPACER ;
    FOREIGN FILL8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 3.680 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 3.680 3.940 ;
        END
    END VDD
END FILL8

MACRO FILL4
    CLASS CORE SPACER ;
    FOREIGN FILL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 1.840 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 1.840 3.940 ;
        END
    END VDD
END FILL4

MACRO FILL2
    CLASS CORE SPACER ;
    FOREIGN FILL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 0.920 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 0.920 3.940 ;
        END
    END VDD
END FILL2

MACRO FILL1
    CLASS CORE SPACER ;
    FOREIGN FILL1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.460 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 0.460 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 0.460 3.940 ;
        END
    END VDD
END FILL1

MACRO ANTENNA
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.330 0.875 0.590 2.385 ;
        RECT  0.125 0.875 0.330 1.185 ;
        END
        ANTENNADIFFAREA     1.4270 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 0.920 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 0.920 3.940 ;
        END
    END VDD
END ANTENNA

MACRO TIELO
    CLASS CORE ;
    FOREIGN TIELO 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 1.105 0.795 1.580 ;
        RECT  0.585 1.035 0.785 1.580 ;
        RECT  0.525 1.035 0.585 1.355 ;
        END
        ANTENNADIFFAREA     0.1428 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 -0.250 0.920 0.250 ;
        RECT  0.125 -0.250 0.725 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 3.440 0.920 3.940 ;
        RECT  0.315 2.700 0.575 3.940 ;
        RECT  0.000 3.440 0.315 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.315 1.760 0.575 2.390 ;
    END
END TIELO

MACRO TIEHI
    CLASS CORE ;
    FOREIGN TIEHI 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 2.110 0.795 2.400 ;
        RECT  0.525 1.955 0.785 2.555 ;
        END
        ANTENNADIFFAREA     0.2176 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 -0.250 0.920 0.250 ;
        RECT  0.385 -0.250 0.645 0.405 ;
        RECT  0.000 -0.250 0.385 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 0.920 3.940 ;
        RECT  0.125 2.875 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.545 1.035 0.645 1.295 ;
        RECT  0.385 1.035 0.545 1.675 ;
        RECT  0.125 1.515 0.385 1.775 ;
    END
END TIEHI

MACRO DLY4X4
    CLASS CORE ;
    FOREIGN DLY4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.105 4.015 1.990 ;
        RECT  3.830 1.005 4.005 1.990 ;
        RECT  3.805 0.880 3.830 1.990 ;
        RECT  3.745 0.880 3.805 1.205 ;
        RECT  3.575 1.790 3.805 1.990 ;
        RECT  3.485 0.605 3.745 1.205 ;
        RECT  3.505 1.790 3.575 2.605 ;
        RECT  3.375 1.790 3.505 3.005 ;
        RECT  3.345 2.335 3.375 3.005 ;
        RECT  3.245 2.405 3.345 3.005 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.295 1.590 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 -0.250 4.140 0.250 ;
        RECT  2.975 -0.250 3.235 1.075 ;
        RECT  0.785 -0.250 2.975 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.255 4.015 3.940 ;
        RECT  2.955 3.440 3.755 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  0.785 3.440 2.695 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.585 3.195 1.845 ;
        RECT  2.935 1.255 3.095 2.220 ;
        RECT  2.155 1.255 2.935 1.415 ;
        RECT  2.155 2.060 2.935 2.220 ;
        RECT  2.275 1.595 2.535 1.855 ;
        RECT  1.725 1.645 2.275 1.805 ;
        RECT  1.995 1.035 2.155 1.415 ;
        RECT  1.995 2.060 2.155 2.770 ;
        RECT  1.895 1.035 1.995 1.295 ;
        RECT  1.895 2.510 1.995 2.770 ;
        RECT  1.715 0.525 1.755 0.785 ;
        RECT  1.715 1.645 1.725 2.260 ;
        RECT  1.555 0.525 1.715 2.260 ;
        RECT  1.495 0.525 1.555 0.785 ;
        RECT  1.465 2.000 1.555 2.260 ;
        RECT  1.135 1.495 1.235 1.755 ;
        RECT  0.975 1.245 1.135 2.330 ;
        RECT  0.385 1.245 0.975 1.405 ;
        RECT  0.385 2.170 0.975 2.330 ;
        RECT  0.125 1.035 0.385 1.405 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END DLY4X4

MACRO DLY3X4
    CLASS CORE ;
    FOREIGN DLY3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.105 4.015 1.990 ;
        RECT  3.830 1.005 4.005 1.990 ;
        RECT  3.805 0.880 3.830 1.990 ;
        RECT  3.745 0.880 3.805 1.205 ;
        RECT  3.575 1.790 3.805 1.990 ;
        RECT  3.485 0.605 3.745 1.205 ;
        RECT  3.505 1.790 3.575 2.605 ;
        RECT  3.375 1.790 3.505 3.005 ;
        RECT  3.345 2.335 3.375 3.005 ;
        RECT  3.245 2.405 3.345 3.005 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.295 1.590 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 -0.250 4.140 0.250 ;
        RECT  2.975 -0.250 3.235 1.075 ;
        RECT  0.785 -0.250 2.975 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.255 4.015 3.940 ;
        RECT  2.955 3.440 3.755 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  0.785 3.440 2.695 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.585 3.195 1.845 ;
        RECT  2.935 1.255 3.095 2.220 ;
        RECT  2.155 1.255 2.935 1.415 ;
        RECT  2.155 2.060 2.935 2.220 ;
        RECT  2.275 1.595 2.535 1.855 ;
        RECT  1.725 1.645 2.275 1.805 ;
        RECT  1.995 1.035 2.155 1.415 ;
        RECT  1.995 2.060 2.155 2.770 ;
        RECT  1.895 1.035 1.995 1.295 ;
        RECT  1.895 2.510 1.995 2.770 ;
        RECT  1.715 0.525 1.755 0.785 ;
        RECT  1.715 1.645 1.725 2.260 ;
        RECT  1.555 0.525 1.715 2.260 ;
        RECT  1.495 0.525 1.555 0.785 ;
        RECT  1.465 2.000 1.555 2.260 ;
        RECT  1.135 1.495 1.235 1.755 ;
        RECT  0.975 1.245 1.135 2.330 ;
        RECT  0.385 1.245 0.975 1.405 ;
        RECT  0.385 2.170 0.975 2.330 ;
        RECT  0.125 1.035 0.385 1.405 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END DLY3X4

MACRO DLY2X4
    CLASS CORE ;
    FOREIGN DLY2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.105 4.015 1.990 ;
        RECT  3.830 1.005 4.005 1.990 ;
        RECT  3.805 0.880 3.830 1.990 ;
        RECT  3.745 0.880 3.805 1.205 ;
        RECT  3.575 1.790 3.805 1.990 ;
        RECT  3.485 0.605 3.745 1.205 ;
        RECT  3.505 1.790 3.575 2.605 ;
        RECT  3.375 1.790 3.505 3.005 ;
        RECT  3.345 2.335 3.375 3.005 ;
        RECT  3.245 2.405 3.345 3.005 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.295 1.590 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 -0.250 4.140 0.250 ;
        RECT  2.975 -0.250 3.235 1.075 ;
        RECT  0.785 -0.250 2.975 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.255 4.015 3.940 ;
        RECT  2.955 3.440 3.755 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  0.785 3.440 2.695 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.585 3.195 1.845 ;
        RECT  2.935 1.255 3.095 2.220 ;
        RECT  2.155 1.255 2.935 1.415 ;
        RECT  2.155 2.060 2.935 2.220 ;
        RECT  2.275 1.595 2.535 1.855 ;
        RECT  1.725 1.645 2.275 1.805 ;
        RECT  1.995 1.035 2.155 1.415 ;
        RECT  1.995 2.060 2.155 2.770 ;
        RECT  1.895 1.035 1.995 1.295 ;
        RECT  1.895 2.510 1.995 2.770 ;
        RECT  1.715 0.525 1.755 0.785 ;
        RECT  1.715 1.645 1.725 2.260 ;
        RECT  1.555 0.525 1.715 2.260 ;
        RECT  1.495 0.525 1.555 0.785 ;
        RECT  1.465 2.000 1.555 2.260 ;
        RECT  1.135 1.495 1.235 1.755 ;
        RECT  0.975 1.245 1.135 2.330 ;
        RECT  0.385 1.245 0.975 1.405 ;
        RECT  0.385 2.170 0.975 2.330 ;
        RECT  0.125 1.035 0.385 1.405 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END DLY2X4

MACRO DLY1X4
    CLASS CORE ;
    FOREIGN DLY1X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.105 4.015 1.990 ;
        RECT  3.830 1.005 4.005 1.990 ;
        RECT  3.805 0.880 3.830 1.990 ;
        RECT  3.745 0.880 3.805 1.205 ;
        RECT  3.575 1.790 3.805 1.990 ;
        RECT  3.485 0.605 3.745 1.205 ;
        RECT  3.505 1.790 3.575 2.605 ;
        RECT  3.375 1.790 3.505 3.005 ;
        RECT  3.345 2.335 3.375 3.005 ;
        RECT  3.245 2.405 3.345 3.005 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.295 1.590 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 -0.250 4.140 0.250 ;
        RECT  2.975 -0.250 3.235 1.075 ;
        RECT  0.785 -0.250 2.975 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.255 4.015 3.940 ;
        RECT  2.955 3.440 3.755 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  0.785 3.440 2.695 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.585 3.195 1.845 ;
        RECT  2.935 1.255 3.095 2.220 ;
        RECT  2.155 1.255 2.935 1.415 ;
        RECT  2.155 2.060 2.935 2.220 ;
        RECT  2.275 1.595 2.535 1.855 ;
        RECT  1.725 1.645 2.275 1.805 ;
        RECT  1.995 1.035 2.155 1.415 ;
        RECT  1.995 2.060 2.155 2.770 ;
        RECT  1.895 1.035 1.995 1.295 ;
        RECT  1.895 2.510 1.995 2.770 ;
        RECT  1.715 0.525 1.755 0.785 ;
        RECT  1.715 1.645 1.725 2.260 ;
        RECT  1.555 0.525 1.715 2.260 ;
        RECT  1.495 0.525 1.555 0.785 ;
        RECT  1.465 2.000 1.555 2.260 ;
        RECT  1.135 1.495 1.235 1.755 ;
        RECT  0.975 1.245 1.135 2.330 ;
        RECT  0.385 1.245 0.975 1.405 ;
        RECT  0.385 2.170 0.975 2.330 ;
        RECT  0.125 1.035 0.385 1.405 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END DLY1X4

MACRO DLY4X1
    CLASS CORE ;
    FOREIGN DLY4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 1.035 3.555 2.555 ;
        RECT  3.370 1.035 3.395 1.355 ;
        RECT  3.370 1.925 3.395 2.555 ;
        RECT  3.295 1.035 3.370 1.295 ;
        RECT  3.295 1.955 3.370 2.555 ;
        END
        ANTENNADIFFAREA     0.3306 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.245 0.795 1.665 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.680 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.785 -0.250 2.835 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.680 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.785 3.440 2.835 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.515 3.195 1.775 ;
        RECT  2.935 1.020 3.095 2.115 ;
        RECT  2.125 1.020 2.935 1.180 ;
        RECT  2.155 1.955 2.935 2.115 ;
        RECT  2.345 1.470 2.605 1.730 ;
        RECT  1.725 1.520 2.345 1.680 ;
        RECT  1.995 1.955 2.155 2.785 ;
        RECT  1.965 0.525 2.125 1.180 ;
        RECT  1.895 2.525 1.995 2.785 ;
        RECT  1.865 0.525 1.965 0.785 ;
        RECT  1.565 1.035 1.725 2.275 ;
        RECT  1.465 1.035 1.565 1.295 ;
        RECT  1.465 2.015 1.565 2.275 ;
        RECT  1.015 1.595 1.265 2.005 ;
        RECT  0.385 1.845 1.015 2.005 ;
        RECT  0.285 0.805 0.385 1.065 ;
        RECT  0.285 1.845 0.385 2.615 ;
        RECT  0.125 0.805 0.285 2.615 ;
    END
END DLY4X1

MACRO DLY3X1
    CLASS CORE ;
    FOREIGN DLY3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 1.035 3.555 2.555 ;
        RECT  3.370 1.035 3.395 1.355 ;
        RECT  3.370 1.925 3.395 2.555 ;
        RECT  3.295 1.035 3.370 1.295 ;
        RECT  3.295 1.955 3.370 2.555 ;
        END
        ANTENNADIFFAREA     0.3306 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.245 0.795 1.665 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.680 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.785 -0.250 2.835 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.680 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.785 3.440 2.835 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.515 3.195 1.775 ;
        RECT  2.935 1.020 3.095 2.115 ;
        RECT  2.125 1.020 2.935 1.180 ;
        RECT  2.155 1.955 2.935 2.115 ;
        RECT  2.345 1.470 2.605 1.730 ;
        RECT  1.725 1.520 2.345 1.680 ;
        RECT  1.995 1.955 2.155 2.785 ;
        RECT  1.965 0.525 2.125 1.180 ;
        RECT  1.895 2.525 1.995 2.785 ;
        RECT  1.865 0.525 1.965 0.785 ;
        RECT  1.565 1.035 1.725 2.275 ;
        RECT  1.465 1.035 1.565 1.295 ;
        RECT  1.465 2.015 1.565 2.275 ;
        RECT  1.015 1.595 1.265 2.005 ;
        RECT  0.385 1.845 1.015 2.005 ;
        RECT  0.285 0.805 0.385 1.065 ;
        RECT  0.285 1.845 0.385 2.615 ;
        RECT  0.125 0.805 0.285 2.615 ;
    END
END DLY3X1

MACRO DLY2X1
    CLASS CORE ;
    FOREIGN DLY2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 1.035 3.555 2.555 ;
        RECT  3.370 1.035 3.395 1.355 ;
        RECT  3.370 1.925 3.395 2.555 ;
        RECT  3.295 1.035 3.370 1.295 ;
        RECT  3.295 1.955 3.370 2.555 ;
        END
        ANTENNADIFFAREA     0.3306 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.245 0.795 1.665 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.680 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.785 -0.250 2.835 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.680 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.785 3.440 2.835 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.515 3.195 1.775 ;
        RECT  2.935 1.020 3.095 2.115 ;
        RECT  2.125 1.020 2.935 1.180 ;
        RECT  2.155 1.955 2.935 2.115 ;
        RECT  2.345 1.470 2.605 1.730 ;
        RECT  1.725 1.520 2.345 1.680 ;
        RECT  1.995 1.955 2.155 2.785 ;
        RECT  1.965 0.525 2.125 1.180 ;
        RECT  1.895 2.525 1.995 2.785 ;
        RECT  1.865 0.525 1.965 0.785 ;
        RECT  1.565 1.035 1.725 2.275 ;
        RECT  1.465 1.035 1.565 1.295 ;
        RECT  1.465 2.015 1.565 2.275 ;
        RECT  1.015 1.595 1.265 2.005 ;
        RECT  0.385 1.845 1.015 2.005 ;
        RECT  0.285 0.805 0.385 1.065 ;
        RECT  0.285 1.845 0.385 2.615 ;
        RECT  0.125 0.805 0.285 2.615 ;
    END
END DLY2X1

MACRO DLY1X1
    CLASS CORE ;
    FOREIGN DLY1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 1.035 3.555 2.555 ;
        RECT  3.370 1.035 3.395 1.355 ;
        RECT  3.370 1.925 3.395 2.555 ;
        RECT  3.295 1.035 3.370 1.295 ;
        RECT  3.295 1.955 3.370 2.555 ;
        END
        ANTENNADIFFAREA     0.3306 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.245 0.795 1.665 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.680 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.785 -0.250 2.835 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.680 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.785 3.440 2.835 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.515 3.195 1.775 ;
        RECT  2.935 1.020 3.095 2.115 ;
        RECT  2.125 1.020 2.935 1.180 ;
        RECT  2.155 1.955 2.935 2.115 ;
        RECT  2.345 1.470 2.605 1.730 ;
        RECT  1.725 1.520 2.345 1.680 ;
        RECT  1.995 1.955 2.155 2.785 ;
        RECT  1.965 0.525 2.125 1.180 ;
        RECT  1.895 2.525 1.995 2.785 ;
        RECT  1.865 0.525 1.965 0.785 ;
        RECT  1.565 1.035 1.725 2.275 ;
        RECT  1.465 1.035 1.565 1.295 ;
        RECT  1.465 2.015 1.565 2.275 ;
        RECT  1.015 1.595 1.265 2.005 ;
        RECT  0.385 1.845 1.015 2.005 ;
        RECT  0.285 0.805 0.385 1.065 ;
        RECT  0.285 1.845 0.385 2.615 ;
        RECT  0.125 0.805 0.285 2.615 ;
    END
END DLY1X1

MACRO RFRDX4
    CLASS CORE ;
    FOREIGN RFRDX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 0.880 2.635 1.355 ;
        RECT  2.450 0.605 2.575 1.480 ;
        RECT  2.415 0.605 2.450 1.580 ;
        RECT  2.315 0.605 2.415 0.865 ;
        RECT  2.325 1.320 2.415 1.580 ;
        RECT  2.165 1.320 2.325 2.215 ;
        RECT  1.335 1.320 2.165 1.480 ;
        RECT  2.065 1.955 2.165 2.215 ;
        RECT  1.075 1.320 1.335 1.665 ;
        END
        ANTENNAGATEAREA     0.5512 ;
        ANTENNADIFFAREA     0.2715 ;
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.625 1.660 1.885 2.050 ;
        RECT  0.900 1.850 1.625 2.050 ;
        RECT  0.895 0.540 0.900 1.140 ;
        RECT  0.895 1.850 0.900 2.895 ;
        RECT  0.640 0.540 0.895 2.895 ;
        RECT  0.585 0.695 0.640 2.585 ;
        END
        ANTENNAGATEAREA     0.1860 ;
        ANTENNADIFFAREA     0.8268 ;
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 -0.250 2.760 0.250 ;
        RECT  1.185 -0.250 1.445 1.140 ;
        RECT  0.385 -0.250 1.185 0.250 ;
        RECT  0.125 -0.250 0.385 1.140 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 3.440 2.760 3.940 ;
        RECT  1.185 2.385 1.445 3.940 ;
        RECT  0.385 3.440 1.185 3.940 ;
        RECT  0.125 2.215 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END RFRDX4

MACRO RFRDX2
    CLASS CORE ;
    FOREIGN RFRDX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 0.605 2.175 1.295 ;
        RECT  1.915 0.605 1.965 0.865 ;
        RECT  1.800 1.130 1.965 1.295 ;
        RECT  1.640 1.130 1.800 2.215 ;
        RECT  0.775 1.320 1.640 1.480 ;
        RECT  1.540 1.955 1.640 2.215 ;
        RECT  0.610 1.320 0.775 1.690 ;
        RECT  0.515 1.430 0.610 1.690 ;
        END
        ANTENNAGATEAREA     0.2756 ;
        ANTENNADIFFAREA     0.3208 ;
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.100 1.660 1.360 2.030 ;
        RECT  0.385 1.870 1.100 2.030 ;
        RECT  0.335 0.625 0.385 1.225 ;
        RECT  0.335 1.870 0.385 3.045 ;
        RECT  0.125 0.625 0.335 3.045 ;
        END
        ANTENNAGATEAREA     0.1860 ;
        ANTENNADIFFAREA     0.7314 ;
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.930 -0.250 2.300 0.250 ;
        RECT  0.670 -0.250 0.930 1.140 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.930 3.440 2.300 3.940 ;
        RECT  0.670 2.215 0.930 3.940 ;
        RECT  0.000 3.440 0.670 3.940 ;
        END
    END VDD
END RFRDX2

MACRO RFRDX1
    CLASS CORE ;
    FOREIGN RFRDX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 0.605 2.175 1.170 ;
        RECT  1.810 0.880 1.915 1.170 ;
        RECT  1.650 0.880 1.810 2.295 ;
        RECT  1.505 1.105 1.650 1.480 ;
        RECT  1.550 2.035 1.650 2.295 ;
        RECT  0.775 1.320 1.505 1.480 ;
        RECT  0.610 1.320 0.775 1.690 ;
        RECT  0.515 1.430 0.610 1.690 ;
        END
        ANTENNAGATEAREA     0.1378 ;
        ANTENNADIFFAREA     0.3209 ;
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.110 1.665 1.370 2.035 ;
        RECT  0.385 1.875 1.110 2.035 ;
        RECT  0.335 0.990 0.385 1.250 ;
        RECT  0.335 1.875 0.385 2.555 ;
        RECT  0.125 0.990 0.335 2.555 ;
        END
        ANTENNAGATEAREA     0.1860 ;
        ANTENNADIFFAREA     0.3657 ;
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.930 -0.250 2.300 0.250 ;
        RECT  0.670 -0.250 0.930 1.140 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.930 3.440 2.300 3.940 ;
        RECT  0.670 2.215 0.930 3.940 ;
        RECT  0.000 3.440 0.670 3.940 ;
        END
    END VDD
END RFRDX1

MACRO RF2R1WX1
    CLASS CORE ;
    FOREIGN RF2R1WX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN WW
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.930 2.635 3.220 ;
        RECT  2.325 2.930 2.425 3.150 ;
        RECT  2.065 2.890 2.325 3.150 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.320 1.275 0.335 1.580 ;
        RECT  0.100 1.275 0.320 1.845 ;
        END
        ANTENNAGATEAREA     0.1807 ;
    END WB
    PIN R2W
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.525 1.430 6.785 1.990 ;
        END
        ANTENNAGATEAREA     0.1716 ;
    END R2W
    PIN R2B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 2.935 6.045 3.195 ;
        RECT  5.855 1.030 5.995 1.290 ;
        RECT  5.685 0.880 5.855 3.195 ;
        RECT  5.645 0.880 5.685 2.995 ;
        END
        ANTENNADIFFAREA     0.5490 ;
    END R2B
    PIN R1W
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.680 1.425 4.935 2.005 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END R1W
    PIN R1B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  4.055 2.935 4.205 3.195 ;
        RECT  4.055 1.035 4.155 1.295 ;
        RECT  3.895 1.035 4.055 3.195 ;
        RECT  3.805 1.700 3.895 2.995 ;
        END
        ANTENNADIFFAREA     0.5536 ;
    END R1B
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.465 -0.250 6.900 0.250 ;
        RECT  6.205 -0.250 6.465 0.575 ;
        RECT  5.055 -0.250 6.205 0.250 ;
        RECT  4.795 -0.250 5.055 0.405 ;
        RECT  3.335 -0.250 4.795 0.250 ;
        RECT  3.175 -0.250 3.335 0.970 ;
        RECT  1.895 -0.250 3.175 0.250 ;
        RECT  1.635 -0.250 1.895 0.755 ;
        RECT  0.385 -0.250 1.635 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 3.440 6.900 3.940 ;
        RECT  6.305 2.895 6.565 3.940 ;
        RECT  5.000 3.440 6.305 3.940 ;
        RECT  5.000 2.860 5.170 3.120 ;
        RECT  4.740 2.860 5.000 3.940 ;
        RECT  4.570 2.860 4.740 3.120 ;
        RECT  3.370 3.440 4.740 3.940 ;
        RECT  3.110 2.390 3.370 3.940 ;
        RECT  1.885 3.440 3.110 3.940 ;
        RECT  1.625 2.690 1.885 3.940 ;
        RECT  0.385 3.440 1.625 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.345 1.025 6.565 1.185 ;
        RECT  6.345 2.265 6.565 2.525 ;
        RECT  6.305 1.025 6.345 2.525 ;
        RECT  6.185 1.025 6.305 2.475 ;
        RECT  6.180 1.745 6.185 2.475 ;
        RECT  6.045 1.745 6.180 2.005 ;
        RECT  5.275 1.400 5.395 1.660 ;
        RECT  5.115 0.685 5.275 1.660 ;
        RECT  3.715 0.685 5.115 0.845 ;
        RECT  4.495 1.085 4.715 1.245 ;
        RECT  4.455 2.275 4.715 2.535 ;
        RECT  4.400 1.085 4.495 1.650 ;
        RECT  4.415 2.275 4.455 2.435 ;
        RECT  4.400 1.905 4.415 2.435 ;
        RECT  4.335 1.085 4.400 2.435 ;
        RECT  4.240 1.490 4.335 2.435 ;
        RECT  3.555 0.685 3.715 1.435 ;
        RECT  3.530 1.275 3.555 1.435 ;
        RECT  3.410 1.275 3.530 1.760 ;
        RECT  3.250 1.275 3.410 2.180 ;
        RECT  2.855 1.275 3.250 1.435 ;
        RECT  2.860 2.020 3.250 2.180 ;
        RECT  2.070 1.615 3.015 1.775 ;
        RECT  2.700 2.020 2.860 2.750 ;
        RECT  2.595 1.035 2.855 1.435 ;
        RECT  2.600 2.490 2.700 2.750 ;
        RECT  1.730 1.275 2.595 1.435 ;
        RECT  2.240 0.525 2.475 0.785 ;
        RECT  2.250 1.955 2.410 2.510 ;
        RECT  1.440 2.350 2.250 2.510 ;
        RECT  2.215 0.525 2.240 1.095 ;
        RECT  2.080 0.575 2.215 1.095 ;
        RECT  1.390 0.935 2.080 1.095 ;
        RECT  1.910 1.615 2.070 2.170 ;
        RECT  1.100 2.010 1.910 2.170 ;
        RECT  1.570 1.275 1.730 1.830 ;
        RECT  1.280 2.350 1.440 3.040 ;
        RECT  1.230 0.695 1.390 1.095 ;
        RECT  0.925 2.880 1.280 3.040 ;
        RECT  0.675 0.695 1.230 0.855 ;
        RECT  1.050 2.010 1.100 2.700 ;
        RECT  0.890 1.035 1.050 2.700 ;
        RECT  0.665 2.880 0.925 3.140 ;
        RECT  0.840 2.100 0.890 2.700 ;
        RECT  0.660 0.695 0.675 1.920 ;
        RECT  0.660 2.880 0.665 3.040 ;
        RECT  0.515 0.695 0.660 3.040 ;
        RECT  0.500 1.760 0.515 3.040 ;
    END
END RF2R1WX1

MACRO RF1R1WX1
    CLASS CORE ;
    FOREIGN RF1R1WX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN WW
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.520 1.715 2.810 ;
        RECT  1.260 2.550 1.505 2.810 ;
        END
        ANTENNAGATEAREA     0.0975 ;
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.370 1.580 0.400 1.840 ;
        RECT  0.125 1.505 0.370 1.990 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END WB
    PIN RWN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.275 2.110 3.555 2.555 ;
        RECT  3.245 2.140 3.275 2.400 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END RWN
    PIN RW
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 0.945 3.200 1.305 ;
        RECT  2.885 0.880 3.095 1.305 ;
        END
        ANTENNAGATEAREA     0.0507 ;
    END RW
    PIN RB
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  3.295 2.735 3.555 2.995 ;
        RECT  3.380 0.505 3.540 1.930 ;
        RECT  3.275 0.505 3.380 0.765 ;
        RECT  3.060 1.770 3.380 1.930 ;
        RECT  3.060 2.735 3.295 2.895 ;
        RECT  2.900 1.770 3.060 2.895 ;
        RECT  2.425 2.520 2.900 2.810 ;
        END
        ANTENNADIFFAREA     0.3984 ;
    END RB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 -0.250 3.680 0.250 ;
        RECT  2.310 -0.250 2.570 0.795 ;
        RECT  0.390 -0.250 2.310 0.250 ;
        RECT  0.130 -0.250 0.390 0.795 ;
        RECT  0.000 -0.250 0.130 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.695 3.440 3.680 3.940 ;
        RECT  2.435 3.285 2.695 3.940 ;
        RECT  1.845 3.440 2.435 3.940 ;
        RECT  1.585 3.285 1.845 3.940 ;
        RECT  0.390 3.440 1.585 3.940 ;
        RECT  0.130 2.885 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.630 1.460 2.720 1.720 ;
        RECT  2.490 1.170 2.630 2.270 ;
        RECT  2.470 1.090 2.490 2.270 ;
        RECT  2.230 1.090 2.470 1.350 ;
        RECT  2.290 2.010 2.470 2.270 ;
        RECT  2.100 1.570 2.290 1.830 ;
        RECT  1.760 1.190 2.230 1.350 ;
        RECT  1.940 1.570 2.100 2.005 ;
        RECT  1.080 1.845 1.940 2.005 ;
        RECT  1.600 1.190 1.760 1.665 ;
        RECT  1.240 0.490 1.500 0.765 ;
        RECT  0.930 2.990 1.300 3.150 ;
        RECT  0.870 0.505 1.240 0.765 ;
        RECT  0.920 1.015 1.080 2.270 ;
        RECT  0.770 2.685 0.930 3.150 ;
        RECT  0.740 0.605 0.870 0.765 ;
        RECT  0.740 2.685 0.770 2.945 ;
        RECT  0.670 0.605 0.740 2.945 ;
        RECT  0.580 0.605 0.670 2.845 ;
    END
END RF1R1WX1

MACRO TLATNSRX4
    CLASS CORE ;
    FOREIGN TLATNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 1.580 0.665 1.840 ;
        RECT  0.335 1.680 0.405 1.840 ;
        RECT  0.125 1.680 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2561 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.305 1.515 6.315 1.990 ;
        RECT  6.145 1.110 6.305 1.990 ;
        RECT  6.105 1.515 6.145 1.990 ;
        END
        ANTENNAGATEAREA     0.4186 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.865 1.105 10.915 2.400 ;
        RECT  10.605 0.655 10.865 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 1.700 9.995 2.400 ;
        RECT  9.585 0.655 9.845 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.885 1.370 7.145 1.630 ;
        RECT  6.775 1.370 6.885 1.580 ;
        RECT  6.565 1.290 6.775 1.580 ;
        END
        ANTENNAGATEAREA     0.1443 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.455 4.545 1.615 ;
        RECT  2.475 1.455 2.635 1.990 ;
        RECT  2.425 1.545 2.475 1.990 ;
        RECT  2.350 1.545 2.425 1.805 ;
        END
        ANTENNAGATEAREA     0.4264 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.375 -0.250 11.500 0.250 ;
        RECT  11.115 -0.250 11.375 1.190 ;
        RECT  10.355 -0.250 11.115 0.250 ;
        RECT  10.095 -0.250 10.355 1.205 ;
        RECT  9.305 -0.250 10.095 0.250 ;
        RECT  9.045 -0.250 9.305 0.405 ;
        RECT  8.535 -0.250 9.045 0.250 ;
        RECT  8.275 -0.250 8.535 0.405 ;
        RECT  7.045 -0.250 8.275 0.250 ;
        RECT  6.785 -0.250 7.045 0.405 ;
        RECT  4.345 -0.250 6.785 0.250 ;
        RECT  4.085 -0.250 4.345 0.590 ;
        RECT  1.005 -0.250 4.085 0.250 ;
        RECT  0.745 -0.250 1.005 0.815 ;
        RECT  0.000 -0.250 0.745 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.375 3.440 11.500 3.940 ;
        RECT  11.115 2.935 11.375 3.940 ;
        RECT  10.355 3.440 11.115 3.940 ;
        RECT  10.095 2.935 10.355 3.940 ;
        RECT  9.305 3.440 10.095 3.940 ;
        RECT  9.045 3.285 9.305 3.940 ;
        RECT  8.385 3.440 9.045 3.940 ;
        RECT  8.125 3.285 8.385 3.940 ;
        RECT  7.045 3.440 8.125 3.940 ;
        RECT  6.785 3.285 7.045 3.940 ;
        RECT  4.965 3.440 6.785 3.940 ;
        RECT  4.705 3.285 4.965 3.940 ;
        RECT  2.685 3.440 4.705 3.940 ;
        RECT  2.425 3.285 2.685 3.940 ;
        RECT  0.935 3.440 2.425 3.940 ;
        RECT  0.675 3.285 0.935 3.940 ;
        RECT  0.000 3.440 0.675 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.145 1.570 11.305 2.755 ;
        RECT  11.095 1.570 11.145 1.830 ;
        RECT  8.935 2.595 11.145 2.755 ;
        RECT  8.835 1.035 8.935 2.845 ;
        RECT  8.775 1.035 8.835 3.100 ;
        RECT  8.675 1.035 8.775 1.295 ;
        RECT  8.675 2.245 8.775 3.100 ;
        RECT  6.405 2.940 8.675 3.100 ;
        RECT  8.485 1.640 8.595 1.900 ;
        RECT  8.435 1.640 8.485 2.760 ;
        RECT  8.325 1.740 8.435 2.760 ;
        RECT  1.465 2.600 8.325 2.760 ;
        RECT  7.895 0.435 8.055 2.415 ;
        RECT  7.685 0.435 7.895 0.595 ;
        RECT  5.825 2.255 7.895 2.415 ;
        RECT  7.555 1.030 7.715 2.075 ;
        RECT  7.455 1.030 7.555 1.190 ;
        RECT  7.215 1.915 7.555 2.075 ;
        RECT  7.360 0.930 7.455 1.190 ;
        RECT  7.195 0.770 7.360 1.190 ;
        RECT  5.465 0.770 7.195 0.930 ;
        RECT  5.925 2.940 6.185 3.200 ;
        RECT  4.275 2.945 5.925 3.105 ;
        RECT  5.665 1.110 5.825 2.415 ;
        RECT  3.965 2.255 5.665 2.415 ;
        RECT  5.125 0.430 5.535 0.590 ;
        RECT  5.335 0.770 5.465 1.275 ;
        RECT  5.305 0.770 5.335 1.680 ;
        RECT  5.075 1.115 5.305 1.680 ;
        RECT  4.965 0.430 5.125 0.930 ;
        RECT  2.660 1.115 5.075 1.275 ;
        RECT  3.185 0.770 4.965 0.930 ;
        RECT  4.015 2.945 4.275 3.260 ;
        RECT  1.375 2.945 4.015 3.105 ;
        RECT  3.705 1.795 3.965 2.415 ;
        RECT  1.985 2.255 3.705 2.415 ;
        RECT  2.905 0.735 3.185 0.930 ;
        RECT  1.565 0.770 2.905 0.930 ;
        RECT  1.825 1.265 1.985 2.415 ;
        RECT  1.465 0.590 1.565 1.190 ;
        RECT  1.305 0.590 1.465 2.760 ;
        RECT  1.125 2.945 1.375 3.225 ;
        RECT  1.115 1.135 1.125 3.225 ;
        RECT  0.965 1.135 1.115 3.105 ;
        RECT  0.495 1.135 0.965 1.295 ;
        RECT  0.395 2.945 0.965 3.105 ;
        RECT  0.235 0.695 0.495 1.295 ;
        RECT  0.135 2.170 0.395 3.110 ;
    END
END TLATNSRX4

MACRO TLATNSRX2
    CLASS CORE ;
    FOREIGN TLATNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.840 ;
        RECT  0.125 1.290 0.335 1.840 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.630 1.475 2.635 1.990 ;
        RECT  2.370 1.475 2.630 2.025 ;
        RECT  2.360 1.475 2.370 1.990 ;
        END
        ANTENNAGATEAREA     0.2288 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 0.655 7.695 3.060 ;
        RECT  7.435 0.655 7.535 1.255 ;
        RECT  7.435 2.120 7.535 3.060 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.615 1.515 6.775 2.400 ;
        RECT  6.565 1.035 6.615 2.400 ;
        RECT  6.465 1.035 6.565 2.335 ;
        RECT  6.455 1.035 6.465 2.215 ;
        RECT  6.355 1.035 6.455 1.295 ;
        RECT  6.415 1.955 6.455 2.215 ;
        END
        ANTENNADIFFAREA     0.6022 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.310 4.550 1.840 ;
        RECT  4.265 1.290 4.475 1.840 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.930 1.455 2.175 1.990 ;
        RECT  1.885 1.580 1.930 1.840 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.155 -0.250 7.820 0.250 ;
        RECT  6.895 -0.250 7.155 0.405 ;
        RECT  5.580 -0.250 6.895 0.250 ;
        RECT  5.320 -0.250 5.580 0.405 ;
        RECT  4.500 -0.250 5.320 0.250 ;
        RECT  4.240 -0.250 4.500 0.405 ;
        RECT  2.065 -0.250 4.240 0.250 ;
        RECT  1.805 -0.250 2.065 0.405 ;
        RECT  0.385 -0.250 1.805 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 3.440 7.820 3.940 ;
        RECT  6.925 2.935 7.185 3.940 ;
        RECT  6.175 3.440 6.925 3.940 ;
        RECT  5.915 3.285 6.175 3.940 ;
        RECT  2.345 3.440 5.915 3.940 ;
        RECT  2.085 3.285 2.345 3.940 ;
        RECT  0.385 3.440 2.085 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.175 1.520 7.355 1.780 ;
        RECT  7.015 0.660 7.175 2.740 ;
        RECT  6.120 0.660 7.015 0.820 ;
        RECT  6.275 2.580 7.015 2.740 ;
        RECT  6.110 2.580 6.275 2.955 ;
        RECT  5.860 0.525 6.120 0.820 ;
        RECT  6.015 2.695 6.110 2.955 ;
        RECT  5.730 2.795 6.015 2.955 ;
        RECT  5.810 1.445 5.980 1.705 ;
        RECT  5.720 1.445 5.810 2.565 ;
        RECT  5.570 2.795 5.730 3.215 ;
        RECT  5.650 1.545 5.720 2.565 ;
        RECT  5.390 2.405 5.650 2.565 ;
        RECT  4.220 3.055 5.570 3.215 ;
        RECT  5.310 0.585 5.470 1.975 ;
        RECT  5.230 2.405 5.390 2.875 ;
        RECT  5.010 0.585 5.310 0.745 ;
        RECT  5.280 1.815 5.310 1.975 ;
        RECT  5.120 1.815 5.280 2.075 ;
        RECT  4.560 2.715 5.230 2.875 ;
        RECT  4.930 1.475 5.130 1.635 ;
        RECT  4.900 2.375 5.050 2.535 ;
        RECT  4.750 0.435 5.010 0.745 ;
        RECT  4.900 0.945 4.930 1.635 ;
        RECT  4.740 0.945 4.900 2.535 ;
        RECT  3.625 0.585 4.750 0.745 ;
        RECT  4.085 0.945 4.740 1.105 ;
        RECT  4.400 2.555 4.560 2.875 ;
        RECT  3.230 2.555 4.400 2.715 ;
        RECT  4.060 2.895 4.220 3.215 ;
        RECT  3.925 0.945 4.085 1.885 ;
        RECT  3.480 1.725 3.925 1.885 ;
        RECT  3.500 0.585 3.625 1.355 ;
        RECT  3.285 2.945 3.545 3.245 ;
        RECT  3.465 0.585 3.500 1.455 ;
        RECT  3.220 1.675 3.480 1.935 ;
        RECT  3.240 1.195 3.465 1.455 ;
        RECT  0.880 2.945 3.285 3.105 ;
        RECT  2.980 0.695 3.240 0.975 ;
        RECT  2.975 1.195 3.240 1.355 ;
        RECT  3.020 2.555 3.230 2.755 ;
        RECT  1.075 2.595 3.020 2.755 ;
        RECT  1.660 0.815 2.980 0.975 ;
        RECT  2.815 1.195 2.975 2.375 ;
        RECT  1.415 2.215 2.815 2.375 ;
        RECT  1.400 0.815 1.660 1.075 ;
        RECT  0.735 0.460 1.495 0.620 ;
        RECT  1.255 1.265 1.415 2.375 ;
        RECT  1.075 0.915 1.400 1.075 ;
        RECT  0.915 0.915 1.075 2.755 ;
        RECT  0.735 2.945 0.880 3.215 ;
        RECT  0.575 0.460 0.735 3.215 ;
    END
END TLATNSRX2

MACRO TLATNSRX1
    CLASS CORE ;
    FOREIGN TLATNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.840 ;
        RECT  0.125 1.290 0.335 1.840 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 1.990 ;
        RECT  2.225 1.675 2.360 1.935 ;
        END
        ANTENNAGATEAREA     0.1391 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.655 0.880 6.775 2.330 ;
        RECT  6.615 0.845 6.655 2.330 ;
        RECT  6.565 0.845 6.615 1.170 ;
        RECT  6.565 1.925 6.615 2.330 ;
        RECT  6.395 0.845 6.565 1.105 ;
        RECT  6.215 2.170 6.565 2.330 ;
        RECT  6.055 2.170 6.215 2.430 ;
        END
        ANTENNADIFFAREA     0.3459 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.870 1.700 6.315 1.990 ;
        RECT  5.975 2.710 6.235 2.970 ;
        RECT  5.870 2.710 5.975 2.870 ;
        RECT  5.710 1.035 5.870 2.870 ;
        END
        ANTENNADIFFAREA     0.3276 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.470 4.325 1.730 ;
        RECT  3.825 1.470 4.015 1.990 ;
        RECT  3.805 1.700 3.825 1.990 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 1.600 2.005 1.860 ;
        RECT  1.745 1.420 1.905 1.860 ;
        RECT  1.715 1.420 1.745 1.580 ;
        RECT  1.505 1.290 1.715 1.580 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.575 -0.250 6.900 0.250 ;
        RECT  6.315 -0.250 6.575 0.405 ;
        RECT  5.295 -0.250 6.315 0.250 ;
        RECT  5.035 -0.250 5.295 0.405 ;
        RECT  4.125 -0.250 5.035 0.250 ;
        RECT  3.865 -0.250 4.125 0.405 ;
        RECT  1.915 -0.250 3.865 0.250 ;
        RECT  1.655 -0.250 1.915 0.405 ;
        RECT  0.385 -0.250 1.655 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.840 6.775 3.940 ;
        RECT  5.610 3.440 6.515 3.940 ;
        RECT  5.350 3.080 5.610 3.940 ;
        RECT  4.480 3.440 5.350 3.940 ;
        RECT  4.220 3.285 4.480 3.940 ;
        RECT  2.385 3.440 4.220 3.940 ;
        RECT  2.125 3.285 2.385 3.940 ;
        RECT  0.385 3.440 2.125 3.940 ;
        RECT  0.125 2.870 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.210 1.360 6.435 1.520 ;
        RECT  6.050 0.590 6.210 1.520 ;
        RECT  5.890 0.590 6.050 0.750 ;
        RECT  5.630 0.465 5.890 0.750 ;
        RECT  5.490 0.590 5.630 0.750 ;
        RECT  5.490 1.600 5.530 2.900 ;
        RECT  5.370 0.590 5.490 2.900 ;
        RECT  5.330 0.590 5.370 1.760 ;
        RECT  4.990 2.740 5.370 2.900 ;
        RECT  5.145 1.955 5.190 2.215 ;
        RECT  4.985 0.690 5.145 2.215 ;
        RECT  4.300 2.400 5.040 2.560 ;
        RECT  4.725 2.740 4.990 3.105 ;
        RECT  4.725 0.690 4.985 0.850 ;
        RECT  4.705 1.080 4.805 2.215 ;
        RECT  4.465 0.490 4.725 0.850 ;
        RECT  4.040 2.945 4.725 3.105 ;
        RECT  4.645 1.030 4.705 2.215 ;
        RECT  4.445 1.030 4.645 1.290 ;
        RECT  4.470 1.955 4.645 2.215 ;
        RECT  3.285 0.690 4.465 0.850 ;
        RECT  3.625 1.130 4.445 1.290 ;
        RECT  4.140 2.400 4.300 2.745 ;
        RECT  1.215 2.585 4.140 2.745 ;
        RECT  3.880 2.945 4.040 3.255 ;
        RECT  3.485 1.130 3.625 2.000 ;
        RECT  3.465 1.130 3.485 2.100 ;
        RECT  3.225 1.840 3.465 2.100 ;
        RECT  3.125 0.690 3.285 1.625 ;
        RECT  3.015 1.410 3.125 1.625 ;
        RECT  2.975 1.465 3.015 1.625 ;
        RECT  2.815 1.465 2.975 2.335 ;
        RECT  2.785 0.950 2.945 1.225 ;
        RECT  2.665 2.945 2.925 3.255 ;
        RECT  1.475 2.175 2.815 2.335 ;
        RECT  1.325 0.950 2.785 1.110 ;
        RECT  0.765 2.945 2.665 3.105 ;
        RECT  1.215 0.510 1.475 0.770 ;
        RECT  1.315 1.760 1.475 2.335 ;
        RECT  1.105 0.950 1.325 1.270 ;
        RECT  0.765 0.610 1.215 0.770 ;
        RECT  1.105 2.535 1.215 2.745 ;
        RECT  0.945 0.950 1.105 2.745 ;
        RECT  0.605 0.610 0.765 3.105 ;
        RECT  0.575 2.745 0.605 3.005 ;
    END
END TLATNSRX1

MACRO TLATNSRXL
    CLASS CORE ;
    FOREIGN TLATNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.850 ;
        RECT  0.125 1.290 0.335 1.850 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 1.990 ;
        RECT  2.225 1.765 2.360 1.925 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 0.880 6.775 2.175 ;
        RECT  6.565 0.865 6.725 2.330 ;
        RECT  6.215 2.170 6.565 2.330 ;
        RECT  6.055 2.170 6.215 2.430 ;
        END
        ANTENNADIFFAREA     0.2585 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.870 1.700 6.315 1.990 ;
        RECT  5.975 2.730 6.235 3.010 ;
        RECT  5.870 1.020 6.030 1.280 ;
        RECT  5.870 2.730 5.975 2.890 ;
        RECT  5.710 1.020 5.870 2.890 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.470 4.375 1.730 ;
        RECT  3.805 1.290 4.015 1.730 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.175 1.580 ;
        RECT  1.925 1.420 1.965 1.580 ;
        RECT  1.765 1.420 1.925 1.965 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.575 -0.250 6.900 0.250 ;
        RECT  6.315 -0.250 6.575 0.405 ;
        RECT  5.295 -0.250 6.315 0.250 ;
        RECT  5.035 -0.250 5.295 0.405 ;
        RECT  4.125 -0.250 5.035 0.250 ;
        RECT  3.865 -0.250 4.125 0.405 ;
        RECT  1.915 -0.250 3.865 0.250 ;
        RECT  1.655 -0.250 1.915 0.405 ;
        RECT  0.385 -0.250 1.655 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.840 6.775 3.940 ;
        RECT  5.610 3.440 6.515 3.940 ;
        RECT  5.350 3.070 5.610 3.940 ;
        RECT  4.480 3.440 5.350 3.940 ;
        RECT  4.220 3.285 4.480 3.940 ;
        RECT  2.235 3.440 4.220 3.940 ;
        RECT  1.975 3.285 2.235 3.940 ;
        RECT  0.385 3.440 1.975 3.940 ;
        RECT  0.125 2.555 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.225 0.610 6.385 1.495 ;
        RECT  6.030 0.610 6.225 0.770 ;
        RECT  5.770 0.510 6.030 0.770 ;
        RECT  5.530 0.610 5.770 0.770 ;
        RECT  5.370 0.610 5.530 2.890 ;
        RECT  4.990 2.730 5.370 2.890 ;
        RECT  5.030 0.690 5.190 2.215 ;
        RECT  4.725 0.690 5.030 0.850 ;
        RECT  4.725 2.730 4.990 3.105 ;
        RECT  4.300 2.390 4.850 2.550 ;
        RECT  4.645 1.030 4.805 2.165 ;
        RECT  4.465 0.520 4.725 0.850 ;
        RECT  4.040 2.945 4.725 3.105 ;
        RECT  4.445 1.030 4.645 1.290 ;
        RECT  3.415 2.005 4.645 2.165 ;
        RECT  3.505 0.690 4.465 0.850 ;
        RECT  4.140 2.390 4.300 2.745 ;
        RECT  1.215 2.585 4.140 2.745 ;
        RECT  3.880 2.945 4.040 3.255 ;
        RECT  3.345 0.690 3.505 1.570 ;
        RECT  3.155 1.840 3.415 2.165 ;
        RECT  2.975 1.410 3.345 1.570 ;
        RECT  2.765 0.950 3.025 1.225 ;
        RECT  2.815 1.410 2.975 2.335 ;
        RECT  2.665 2.945 2.925 3.255 ;
        RECT  1.445 2.175 2.815 2.335 ;
        RECT  1.325 0.950 2.765 1.110 ;
        RECT  0.765 2.945 2.665 3.105 ;
        RECT  0.765 0.610 1.535 0.770 ;
        RECT  1.285 1.705 1.445 2.335 ;
        RECT  1.105 0.950 1.325 1.250 ;
        RECT  1.105 2.535 1.215 2.745 ;
        RECT  0.945 0.950 1.105 2.745 ;
        RECT  0.605 0.610 0.765 3.105 ;
        RECT  0.600 2.685 0.605 2.945 ;
    END
END TLATNSRXL

MACRO TLATNX4
    CLASS CORE ;
    FOREIGN TLATNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 1.105 6.775 1.990 ;
        RECT  6.465 0.695 6.725 2.220 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.705 1.290 5.855 1.990 ;
        RECT  5.445 0.695 5.705 2.220 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 0.880 0.370 1.895 ;
        RECT  0.110 1.515 0.125 1.895 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 1.485 1.835 1.990 ;
        RECT  1.505 1.700 1.575 1.990 ;
        END
        ANTENNAGATEAREA     0.4628 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 -0.250 7.360 0.250 ;
        RECT  6.975 -0.250 7.235 1.095 ;
        RECT  6.215 -0.250 6.975 0.250 ;
        RECT  5.955 -0.250 6.215 1.095 ;
        RECT  5.190 -0.250 5.955 0.250 ;
        RECT  4.930 -0.250 5.190 1.095 ;
        RECT  3.485 -0.250 4.930 0.250 ;
        RECT  3.225 -0.250 3.485 0.405 ;
        RECT  1.695 -0.250 3.225 0.250 ;
        RECT  1.435 -0.250 1.695 0.735 ;
        RECT  0.385 -0.250 1.435 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 3.440 7.360 3.940 ;
        RECT  6.975 2.940 7.235 3.940 ;
        RECT  6.215 3.440 6.975 3.940 ;
        RECT  5.955 2.940 6.215 3.940 ;
        RECT  5.165 3.440 5.955 3.940 ;
        RECT  4.905 3.285 5.165 3.940 ;
        RECT  3.220 3.440 4.905 3.940 ;
        RECT  3.060 2.955 3.220 3.940 ;
        RECT  1.580 3.440 3.060 3.940 ;
        RECT  1.320 2.955 1.580 3.940 ;
        RECT  0.385 3.440 1.320 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.150 1.580 7.250 1.840 ;
        RECT  6.990 1.580 7.150 2.760 ;
        RECT  5.225 2.600 6.990 2.760 ;
        RECT  5.065 1.280 5.225 2.760 ;
        RECT  4.725 1.280 5.065 1.440 ;
        RECT  4.725 2.600 5.065 2.760 ;
        RECT  4.355 1.795 4.885 2.055 ;
        RECT  4.610 0.655 4.725 1.440 ;
        RECT  4.465 2.600 4.725 2.910 ;
        RECT  4.565 0.555 4.610 1.440 ;
        RECT  4.350 0.555 4.565 0.815 ;
        RECT  3.590 2.750 4.465 2.910 ;
        RECT  4.270 1.115 4.355 2.055 ;
        RECT  3.985 0.655 4.350 0.815 ;
        RECT  4.195 1.115 4.270 2.420 ;
        RECT  3.475 1.115 4.195 1.275 ;
        RECT  4.110 1.895 4.195 2.420 ;
        RECT  3.175 2.260 4.110 2.420 ;
        RECT  3.855 1.455 4.015 1.715 ;
        RECT  3.725 0.475 3.985 0.815 ;
        RECT  3.135 1.455 3.855 1.615 ;
        RECT  3.430 2.750 3.590 3.120 ;
        RECT  2.795 1.815 3.585 1.975 ;
        RECT  3.315 0.795 3.475 1.275 ;
        RECT  2.585 0.795 3.315 0.955 ;
        RECT  3.015 2.260 3.175 2.775 ;
        RECT  2.975 1.145 3.135 1.615 ;
        RECT  2.435 2.615 3.015 2.775 ;
        RECT  2.215 1.145 2.975 1.305 ;
        RECT  2.695 1.485 2.795 1.975 ;
        RECT  2.535 1.485 2.695 2.410 ;
        RECT  2.325 0.695 2.585 0.955 ;
        RECT  1.995 2.250 2.535 2.410 ;
        RECT  2.175 2.615 2.435 3.215 ;
        RECT  2.215 1.805 2.315 2.065 ;
        RECT  2.055 1.145 2.215 2.065 ;
        RECT  1.265 1.145 2.055 1.305 ;
        RECT  1.835 2.250 1.995 2.740 ;
        RECT  0.785 2.580 1.835 2.740 ;
        RECT  1.185 1.140 1.265 2.400 ;
        RECT  1.105 0.525 1.185 2.400 ;
        RECT  1.025 0.525 1.105 1.305 ;
        RECT  0.925 2.140 1.105 2.400 ;
        RECT  0.925 0.525 1.025 0.785 ;
        RECT  0.710 1.640 0.925 1.900 ;
        RECT  0.710 1.035 0.815 1.295 ;
        RECT  0.710 2.580 0.785 2.910 ;
        RECT  0.550 1.035 0.710 2.910 ;
        RECT  0.525 2.650 0.550 2.910 ;
    END
END TLATNX4

MACRO TLATNX2
    CLASS CORE ;
    FOREIGN TLATNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.390 0.695 5.395 0.945 ;
        RECT  5.390 2.335 5.395 2.995 ;
        RECT  5.230 0.575 5.390 3.045 ;
        RECT  5.130 0.575 5.230 1.175 ;
        RECT  5.130 2.105 5.230 3.045 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 1.515 4.475 1.990 ;
        RECT  4.310 1.515 4.340 2.900 ;
        RECT  4.080 1.035 4.310 2.900 ;
        RECT  4.050 1.035 4.080 1.295 ;
        END
        ANTENNADIFFAREA     0.6988 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.475 0.445 1.735 ;
        RECT  0.335 1.260 0.360 1.735 ;
        RECT  0.125 1.260 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0832 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.680 1.290 1.715 1.580 ;
        RECT  1.395 1.085 1.680 1.600 ;
        END
        ANTENNAGATEAREA     0.2522 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.850 -0.250 5.520 0.250 ;
        RECT  4.590 -0.250 4.850 0.405 ;
        RECT  3.260 -0.250 4.590 0.250 ;
        RECT  3.000 -0.250 3.260 0.925 ;
        RECT  1.465 -0.250 3.000 0.250 ;
        RECT  1.205 -0.250 1.465 0.405 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.850 3.440 5.520 3.940 ;
        RECT  4.590 2.245 4.850 3.940 ;
        RECT  3.220 3.440 4.590 3.940 ;
        RECT  2.960 2.485 3.220 3.940 ;
        RECT  1.360 3.440 2.960 3.940 ;
        RECT  1.100 3.285 1.360 3.940 ;
        RECT  0.385 3.440 1.100 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.950 1.405 5.050 1.665 ;
        RECT  4.790 0.695 4.950 1.665 ;
        RECT  3.800 0.695 4.790 0.855 ;
        RECT  3.705 2.420 3.830 2.680 ;
        RECT  3.705 0.695 3.800 1.005 ;
        RECT  3.545 0.695 3.705 2.680 ;
        RECT  3.540 0.695 3.545 1.005 ;
        RECT  2.960 1.990 3.545 2.250 ;
        RECT  2.780 1.220 3.365 1.480 ;
        RECT  2.620 1.220 2.780 2.755 ;
        RECT  2.315 1.220 2.620 1.380 ;
        RECT  2.230 2.595 2.620 2.755 ;
        RECT  2.315 0.445 2.575 0.745 ;
        RECT  2.280 2.145 2.440 2.410 ;
        RECT  1.215 0.585 2.315 0.745 ;
        RECT  2.155 0.965 2.315 1.380 ;
        RECT  1.715 2.250 2.280 2.410 ;
        RECT  1.970 2.595 2.230 3.195 ;
        RECT  2.055 0.965 2.155 1.225 ;
        RECT  1.895 1.665 2.155 1.945 ;
        RECT  1.215 1.785 1.895 1.945 ;
        RECT  1.555 2.250 1.715 3.105 ;
        RECT  0.380 2.945 1.555 3.105 ;
        RECT  1.055 0.585 1.215 2.765 ;
        RECT  0.895 0.585 1.055 0.785 ;
        RECT  0.560 2.605 1.055 2.765 ;
        RECT  0.635 0.525 0.895 0.785 ;
        RECT  0.815 1.515 0.875 1.840 ;
        RECT  0.655 1.035 0.815 2.330 ;
        RECT  0.555 1.035 0.655 1.295 ;
        RECT  0.525 1.955 0.655 2.330 ;
        RECT  0.380 2.170 0.525 2.330 ;
        RECT  0.220 2.170 0.380 3.105 ;
    END
END TLATNX2

MACRO TLATNX1
    CLASS CORE ;
    FOREIGN TLATNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.025 4.475 2.810 ;
        RECT  4.255 1.025 4.265 1.285 ;
        RECT  4.215 2.305 4.265 2.565 ;
        END
        ANTENNADIFFAREA     0.4535 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.035 0.595 4.075 2.125 ;
        RECT  3.915 0.595 4.035 2.855 ;
        RECT  3.680 0.595 3.915 0.755 ;
        RECT  3.875 1.965 3.915 2.855 ;
        RECT  3.805 2.520 3.875 2.855 ;
        RECT  3.250 2.595 3.805 2.855 ;
        RECT  3.420 0.430 3.680 0.755 ;
        END
        ANTENNADIFFAREA     0.3691 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.475 0.445 1.735 ;
        RECT  0.335 1.260 0.360 1.735 ;
        RECT  0.125 1.260 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.680 1.290 1.715 1.580 ;
        RECT  1.395 1.080 1.680 1.595 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.270 -0.250 4.600 0.250 ;
        RECT  4.010 -0.250 4.270 0.405 ;
        RECT  3.055 -0.250 4.010 0.250 ;
        RECT  2.795 -0.250 3.055 0.405 ;
        RECT  1.475 -0.250 2.795 0.250 ;
        RECT  1.215 -0.250 1.475 0.405 ;
        RECT  0.385 -0.250 1.215 0.250 ;
        RECT  0.125 -0.250 0.385 0.805 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 3.440 4.600 3.940 ;
        RECT  3.620 3.285 3.880 3.940 ;
        RECT  2.925 3.440 3.620 3.940 ;
        RECT  2.665 3.285 2.925 3.940 ;
        RECT  1.325 3.440 2.665 3.940 ;
        RECT  1.065 3.065 1.325 3.940 ;
        RECT  0.385 3.440 1.065 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.635 1.500 3.735 1.760 ;
        RECT  3.475 1.125 3.635 2.295 ;
        RECT  3.375 1.125 3.475 1.385 ;
        RECT  2.985 2.135 3.475 2.295 ;
        RECT  2.645 1.685 3.255 1.945 ;
        RECT  2.825 2.135 2.985 3.075 ;
        RECT  2.375 2.915 2.825 3.075 ;
        RECT  2.485 1.025 2.645 2.435 ;
        RECT  2.255 0.485 2.515 0.745 ;
        RECT  2.285 1.025 2.485 1.185 ;
        RECT  2.065 2.275 2.485 2.435 ;
        RECT  2.025 0.925 2.285 1.185 ;
        RECT  1.215 0.585 2.255 0.745 ;
        RECT  1.805 2.175 2.065 2.435 ;
        RECT  1.215 1.775 1.905 1.935 ;
        RECT  1.055 0.585 1.215 2.555 ;
        RECT  0.895 0.585 1.055 0.785 ;
        RECT  0.745 2.395 1.055 2.555 ;
        RECT  0.635 0.525 0.895 0.785 ;
        RECT  0.815 1.515 0.875 1.840 ;
        RECT  0.655 1.035 0.815 2.215 ;
        RECT  0.585 2.395 0.745 2.815 ;
        RECT  0.555 1.035 0.655 1.295 ;
        RECT  0.525 1.955 0.655 2.215 ;
        RECT  0.485 2.555 0.585 2.815 ;
    END
END TLATNX1

MACRO TLATNXL
    CLASS CORE ;
    FOREIGN TLATNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.025 4.475 2.565 ;
        RECT  4.215 2.305 4.265 2.565 ;
        END
        ANTENNADIFFAREA     0.2827 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 0.625 4.075 2.125 ;
        RECT  3.915 0.625 3.970 2.680 ;
        RECT  3.680 0.625 3.915 0.785 ;
        RECT  3.810 1.965 3.915 2.680 ;
        RECT  3.555 2.520 3.810 2.680 ;
        RECT  3.420 0.525 3.680 0.785 ;
        RECT  3.510 2.520 3.555 2.810 ;
        RECT  3.250 2.520 3.510 2.855 ;
        END
        ANTENNADIFFAREA     0.2340 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.475 0.445 1.735 ;
        RECT  0.125 1.300 0.360 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.670 1.290 1.715 1.580 ;
        RECT  1.395 1.080 1.670 1.595 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.280 -0.250 4.600 0.250 ;
        RECT  4.020 -0.250 4.280 0.405 ;
        RECT  3.095 -0.250 4.020 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  1.465 -0.250 2.835 0.250 ;
        RECT  1.205 -0.250 1.465 0.405 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.805 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 3.440 4.600 3.940 ;
        RECT  3.620 3.285 3.880 3.940 ;
        RECT  3.035 3.440 3.620 3.940 ;
        RECT  2.775 3.285 3.035 3.940 ;
        RECT  1.385 3.440 2.775 3.940 ;
        RECT  1.125 3.285 1.385 3.940 ;
        RECT  0.385 3.440 1.125 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.630 1.500 3.735 1.760 ;
        RECT  3.630 1.035 3.680 1.295 ;
        RECT  3.470 1.035 3.630 2.295 ;
        RECT  3.420 1.035 3.470 1.295 ;
        RECT  2.985 2.135 3.470 2.295 ;
        RECT  2.870 1.685 3.255 1.945 ;
        RECT  2.825 2.135 2.985 3.060 ;
        RECT  2.710 0.735 2.870 1.945 ;
        RECT  2.595 2.900 2.825 3.060 ;
        RECT  2.315 0.735 2.710 0.895 ;
        RECT  2.645 1.785 2.710 1.945 ;
        RECT  2.485 1.785 2.645 2.370 ;
        RECT  2.335 2.900 2.595 3.160 ;
        RECT  2.305 1.080 2.515 1.240 ;
        RECT  2.125 2.210 2.485 2.370 ;
        RECT  2.055 0.635 2.315 0.895 ;
        RECT  2.145 1.080 2.305 2.030 ;
        RECT  1.215 1.870 2.145 2.030 ;
        RECT  1.865 2.210 2.125 2.470 ;
        RECT  1.810 2.900 2.070 3.160 ;
        RECT  0.305 2.945 1.810 3.105 ;
        RECT  1.055 0.590 1.215 2.765 ;
        RECT  0.895 0.590 1.055 0.750 ;
        RECT  0.485 2.605 1.055 2.765 ;
        RECT  0.635 0.430 0.895 0.750 ;
        RECT  0.815 1.515 0.875 1.780 ;
        RECT  0.655 1.035 0.815 2.330 ;
        RECT  0.555 1.035 0.655 1.295 ;
        RECT  0.555 1.960 0.655 2.330 ;
        RECT  0.305 2.170 0.555 2.330 ;
        RECT  0.145 2.170 0.305 3.105 ;
    END
END TLATNXL

MACRO TLATSRX4
    CLASS CORE ;
    FOREIGN TLATSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 1.580 0.665 1.860 ;
        RECT  0.335 1.700 0.405 1.860 ;
        RECT  0.125 1.700 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2561 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.105 1.195 6.405 1.730 ;
        END
        ANTENNAGATEAREA     0.4212 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.855 1.105 10.915 2.400 ;
        RECT  10.595 0.655 10.855 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.835 1.700 9.995 2.400 ;
        RECT  9.575 0.655 9.835 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.855 1.290 7.235 1.665 ;
        END
        ANTENNAGATEAREA     0.1443 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.445 1.445 4.705 1.615 ;
        RECT  2.745 1.445 4.445 1.605 ;
        RECT  2.635 1.445 2.745 1.925 ;
        RECT  2.585 1.445 2.635 1.990 ;
        RECT  2.485 1.535 2.585 1.990 ;
        RECT  2.425 1.700 2.485 1.990 ;
        END
        ANTENNAGATEAREA     0.4264 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.365 -0.250 11.500 0.250 ;
        RECT  11.105 -0.250 11.365 1.190 ;
        RECT  10.345 -0.250 11.105 0.250 ;
        RECT  10.085 -0.250 10.345 1.205 ;
        RECT  9.285 -0.250 10.085 0.250 ;
        RECT  9.025 -0.250 9.285 0.405 ;
        RECT  8.525 -0.250 9.025 0.250 ;
        RECT  8.265 -0.250 8.525 0.405 ;
        RECT  7.145 -0.250 8.265 0.250 ;
        RECT  6.885 -0.250 7.145 0.405 ;
        RECT  4.500 -0.250 6.885 0.250 ;
        RECT  4.240 -0.250 4.500 0.585 ;
        RECT  0.935 -0.250 4.240 0.250 ;
        RECT  0.675 -0.250 0.935 0.945 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.370 3.440 11.500 3.940 ;
        RECT  11.110 2.935 11.370 3.940 ;
        RECT  10.345 3.440 11.110 3.940 ;
        RECT  10.085 2.935 10.345 3.940 ;
        RECT  9.285 3.440 10.085 3.940 ;
        RECT  9.025 3.285 9.285 3.940 ;
        RECT  8.365 3.440 9.025 3.940 ;
        RECT  8.105 3.285 8.365 3.940 ;
        RECT  7.040 3.440 8.105 3.940 ;
        RECT  6.780 3.285 7.040 3.940 ;
        RECT  4.815 3.440 6.780 3.940 ;
        RECT  4.555 3.285 4.815 3.940 ;
        RECT  2.685 3.440 4.555 3.940 ;
        RECT  2.425 3.285 2.685 3.940 ;
        RECT  0.935 3.440 2.425 3.940 ;
        RECT  0.675 3.285 0.935 3.940 ;
        RECT  0.000 3.440 0.675 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.095 1.570 11.255 2.755 ;
        RECT  8.925 2.595 11.095 2.755 ;
        RECT  8.825 1.035 8.925 2.845 ;
        RECT  8.765 1.035 8.825 3.105 ;
        RECT  8.665 1.035 8.765 1.295 ;
        RECT  8.665 2.245 8.765 3.105 ;
        RECT  6.410 2.945 8.665 3.105 ;
        RECT  8.485 1.785 8.585 2.045 ;
        RECT  8.325 1.785 8.485 2.760 ;
        RECT  1.520 2.600 8.325 2.760 ;
        RECT  7.935 0.610 8.085 2.370 ;
        RECT  7.925 0.435 7.935 2.370 ;
        RECT  7.675 0.435 7.925 0.770 ;
        RECT  7.690 2.210 7.925 2.370 ;
        RECT  7.575 1.470 7.745 1.730 ;
        RECT  7.000 0.610 7.675 0.770 ;
        RECT  7.440 0.950 7.575 2.005 ;
        RECT  7.415 0.950 7.440 2.415 ;
        RECT  7.285 0.950 7.415 1.110 ;
        RECT  7.280 1.845 7.415 2.415 ;
        RECT  7.180 2.115 7.280 2.415 ;
        RECT  5.925 2.255 7.180 2.415 ;
        RECT  6.840 0.610 7.000 0.935 ;
        RECT  5.575 0.775 6.840 0.935 ;
        RECT  4.275 2.945 6.190 3.105 ;
        RECT  5.765 1.115 5.925 2.415 ;
        RECT  3.965 2.255 5.765 2.415 ;
        RECT  5.235 0.430 5.705 0.590 ;
        RECT  5.495 0.775 5.575 1.265 ;
        RECT  5.415 0.775 5.495 1.685 ;
        RECT  5.235 1.105 5.415 1.685 ;
        RECT  5.075 0.430 5.235 0.925 ;
        RECT  3.055 1.105 5.235 1.265 ;
        RECT  3.440 0.765 5.075 0.925 ;
        RECT  4.015 2.945 4.275 3.235 ;
        RECT  1.375 2.945 4.015 3.105 ;
        RECT  3.705 1.785 3.965 2.415 ;
        RECT  2.105 2.255 3.705 2.415 ;
        RECT  3.280 0.665 3.440 0.925 ;
        RECT  1.520 0.665 3.280 0.825 ;
        RECT  2.795 1.005 3.055 1.265 ;
        RECT  1.945 1.250 2.105 2.415 ;
        RECT  1.360 0.625 1.520 2.760 ;
        RECT  1.115 2.945 1.375 3.230 ;
        RECT  1.185 0.625 1.360 1.225 ;
        RECT  1.255 2.160 1.360 2.760 ;
        RECT  1.005 1.405 1.180 1.665 ;
        RECT  1.005 2.945 1.115 3.105 ;
        RECT  0.845 1.135 1.005 3.105 ;
        RECT  0.425 1.135 0.845 1.295 ;
        RECT  0.385 2.945 0.845 3.105 ;
        RECT  0.165 0.695 0.425 1.295 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END TLATSRX4

MACRO TLATSRX2
    CLASS CORE ;
    FOREIGN TLATSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.840 ;
        RECT  0.125 1.290 0.335 1.840 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 2.025 ;
        END
        ANTENNAGATEAREA     0.2288 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 0.655 7.695 3.060 ;
        RECT  7.435 0.655 7.535 1.255 ;
        RECT  7.435 2.120 7.535 3.060 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.615 1.515 6.775 2.400 ;
        RECT  6.565 1.035 6.615 2.400 ;
        RECT  6.455 1.035 6.565 2.215 ;
        RECT  6.355 1.035 6.455 1.295 ;
        RECT  6.415 1.955 6.455 2.215 ;
        END
        ANTENNADIFFAREA     0.5833 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.310 4.550 1.840 ;
        RECT  4.265 1.290 4.475 1.840 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 1.290 2.175 1.845 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.155 -0.250 7.820 0.250 ;
        RECT  6.895 -0.250 7.155 0.405 ;
        RECT  5.580 -0.250 6.895 0.250 ;
        RECT  5.320 -0.250 5.580 0.405 ;
        RECT  4.500 -0.250 5.320 0.250 ;
        RECT  4.240 -0.250 4.500 0.405 ;
        RECT  2.065 -0.250 4.240 0.250 ;
        RECT  1.805 -0.250 2.065 0.405 ;
        RECT  0.385 -0.250 1.805 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 3.440 7.820 3.940 ;
        RECT  6.925 2.935 7.185 3.940 ;
        RECT  6.175 3.440 6.925 3.940 ;
        RECT  5.915 3.285 6.175 3.940 ;
        RECT  2.345 3.440 5.915 3.940 ;
        RECT  2.085 3.285 2.345 3.940 ;
        RECT  0.385 3.440 2.085 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.175 1.520 7.355 1.780 ;
        RECT  7.015 0.660 7.175 2.740 ;
        RECT  6.150 0.660 7.015 0.820 ;
        RECT  6.275 2.580 7.015 2.740 ;
        RECT  6.175 2.465 6.275 2.740 ;
        RECT  6.015 2.465 6.175 2.955 ;
        RECT  5.890 0.525 6.150 0.820 ;
        RECT  5.730 2.795 6.015 2.955 ;
        RECT  5.810 1.445 5.980 1.705 ;
        RECT  5.720 1.445 5.810 2.565 ;
        RECT  5.570 2.795 5.730 3.215 ;
        RECT  5.650 1.545 5.720 2.565 ;
        RECT  5.390 2.405 5.650 2.565 ;
        RECT  4.220 3.055 5.570 3.215 ;
        RECT  5.310 0.865 5.470 1.975 ;
        RECT  5.230 2.405 5.390 2.875 ;
        RECT  5.295 0.865 5.310 1.025 ;
        RECT  5.280 1.815 5.310 1.975 ;
        RECT  5.135 0.585 5.295 1.025 ;
        RECT  5.120 1.815 5.280 2.075 ;
        RECT  4.560 2.715 5.230 2.875 ;
        RECT  5.010 0.585 5.135 0.745 ;
        RECT  4.930 1.475 5.130 1.635 ;
        RECT  4.900 2.375 5.050 2.535 ;
        RECT  4.750 0.435 5.010 0.745 ;
        RECT  4.900 0.945 4.930 1.635 ;
        RECT  4.740 0.945 4.900 2.535 ;
        RECT  4.085 0.585 4.750 0.745 ;
        RECT  4.670 0.945 4.740 1.105 ;
        RECT  2.975 2.215 4.740 2.375 ;
        RECT  4.400 2.555 4.560 2.875 ;
        RECT  1.075 2.555 4.400 2.715 ;
        RECT  4.060 2.895 4.220 3.215 ;
        RECT  3.925 0.585 4.085 1.835 ;
        RECT  3.480 1.675 3.925 1.835 ;
        RECT  3.285 2.945 3.545 3.245 ;
        RECT  2.975 1.195 3.500 1.455 ;
        RECT  3.220 1.675 3.480 1.935 ;
        RECT  0.880 2.945 3.285 3.105 ;
        RECT  2.980 0.695 3.240 0.975 ;
        RECT  1.660 0.815 2.980 0.975 ;
        RECT  2.815 1.195 2.975 2.375 ;
        RECT  1.415 2.215 2.815 2.375 ;
        RECT  1.400 0.815 1.660 1.075 ;
        RECT  0.735 0.460 1.495 0.620 ;
        RECT  1.255 1.265 1.415 2.375 ;
        RECT  1.075 0.915 1.400 1.075 ;
        RECT  0.915 0.915 1.075 2.715 ;
        RECT  0.735 2.945 0.880 3.255 ;
        RECT  0.575 0.460 0.735 3.255 ;
    END
END TLATSRX2

MACRO TLATSRX1
    CLASS CORE ;
    FOREIGN TLATSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.840 ;
        RECT  0.125 1.290 0.335 1.840 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 1.990 ;
        RECT  2.225 1.675 2.360 1.935 ;
        END
        ANTENNAGATEAREA     0.1391 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 0.880 6.775 2.180 ;
        RECT  6.565 0.880 6.725 2.330 ;
        RECT  6.395 0.895 6.565 1.055 ;
        RECT  6.215 2.170 6.565 2.330 ;
        RECT  6.055 2.170 6.215 2.430 ;
        END
        ANTENNADIFFAREA     0.3459 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.870 1.700 6.315 1.990 ;
        RECT  6.135 2.950 6.235 3.210 ;
        RECT  5.975 2.730 6.135 3.210 ;
        RECT  5.870 2.730 5.975 2.890 ;
        RECT  5.710 1.035 5.870 2.890 ;
        END
        ANTENNADIFFAREA     0.3276 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.260 1.420 4.325 1.705 ;
        RECT  4.015 1.375 4.260 1.705 ;
        RECT  3.805 1.290 4.015 1.705 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 1.600 2.005 1.860 ;
        RECT  1.745 1.420 1.905 1.860 ;
        RECT  1.715 1.420 1.745 1.580 ;
        RECT  1.505 1.290 1.715 1.580 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.575 -0.250 6.900 0.250 ;
        RECT  6.315 -0.250 6.575 0.405 ;
        RECT  5.295 -0.250 6.315 0.250 ;
        RECT  5.035 -0.250 5.295 0.405 ;
        RECT  4.125 -0.250 5.035 0.250 ;
        RECT  3.865 -0.250 4.125 0.405 ;
        RECT  1.915 -0.250 3.865 0.250 ;
        RECT  1.655 -0.250 1.915 0.405 ;
        RECT  0.385 -0.250 1.655 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.840 6.775 3.940 ;
        RECT  5.695 3.440 6.515 3.940 ;
        RECT  5.435 3.080 5.695 3.940 ;
        RECT  4.470 3.440 5.435 3.940 ;
        RECT  4.210 3.285 4.470 3.940 ;
        RECT  2.380 3.440 4.210 3.940 ;
        RECT  2.120 3.285 2.380 3.940 ;
        RECT  0.385 3.440 2.120 3.940 ;
        RECT  0.125 2.870 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.225 1.260 6.385 1.520 ;
        RECT  6.210 1.260 6.225 1.420 ;
        RECT  6.050 0.590 6.210 1.420 ;
        RECT  5.890 0.590 6.050 0.750 ;
        RECT  5.630 0.465 5.890 0.750 ;
        RECT  5.490 0.590 5.630 0.750 ;
        RECT  5.490 1.600 5.530 2.900 ;
        RECT  5.370 0.590 5.490 2.900 ;
        RECT  5.330 0.590 5.370 1.760 ;
        RECT  5.120 2.740 5.370 2.900 ;
        RECT  5.145 1.955 5.190 2.215 ;
        RECT  4.985 0.700 5.145 2.215 ;
        RECT  4.860 2.740 5.120 3.105 ;
        RECT  4.300 2.400 5.040 2.560 ;
        RECT  4.725 0.700 4.985 0.860 ;
        RECT  4.030 2.945 4.860 3.105 ;
        RECT  4.645 1.080 4.805 2.215 ;
        RECT  4.465 0.520 4.725 0.860 ;
        RECT  4.445 1.080 4.645 1.240 ;
        RECT  4.470 1.955 4.645 2.215 ;
        RECT  3.960 2.055 4.470 2.215 ;
        RECT  3.615 0.700 4.465 0.860 ;
        RECT  4.140 2.400 4.300 2.745 ;
        RECT  1.210 2.585 4.140 2.745 ;
        RECT  3.870 2.945 4.030 3.255 ;
        RECT  3.800 2.055 3.960 2.405 ;
        RECT  2.975 2.245 3.800 2.405 ;
        RECT  3.455 0.700 3.615 2.050 ;
        RECT  3.155 1.890 3.455 2.050 ;
        RECT  2.975 1.410 3.275 1.570 ;
        RECT  2.765 0.950 3.025 1.225 ;
        RECT  2.815 1.410 2.975 2.405 ;
        RECT  2.660 2.945 2.920 3.255 ;
        RECT  1.475 2.175 2.815 2.335 ;
        RECT  1.325 0.950 2.765 1.110 ;
        RECT  0.755 2.945 2.660 3.105 ;
        RECT  1.215 0.510 1.475 0.770 ;
        RECT  1.315 1.760 1.475 2.335 ;
        RECT  1.105 0.950 1.325 1.270 ;
        RECT  0.740 0.610 1.215 0.770 ;
        RECT  1.105 2.515 1.210 2.745 ;
        RECT  0.945 0.950 1.105 2.745 ;
        RECT  0.740 1.035 0.765 1.295 ;
        RECT  0.740 2.795 0.755 3.105 ;
        RECT  0.595 0.610 0.740 3.105 ;
        RECT  0.580 0.610 0.595 3.005 ;
        RECT  0.565 2.745 0.580 3.005 ;
    END
END TLATSRX1

MACRO TLATSRXL
    CLASS CORE ;
    FOREIGN TLATSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.850 ;
        RECT  0.125 1.290 0.335 1.850 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 1.990 ;
        RECT  2.225 1.760 2.360 1.920 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 0.880 6.775 2.175 ;
        RECT  6.565 0.865 6.725 2.330 ;
        RECT  6.215 2.170 6.565 2.330 ;
        RECT  6.055 2.170 6.215 2.430 ;
        END
        ANTENNADIFFAREA     0.2585 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.870 1.700 6.315 1.990 ;
        RECT  5.975 2.730 6.235 3.010 ;
        RECT  5.870 1.020 6.030 1.280 ;
        RECT  5.870 2.730 5.975 2.890 ;
        RECT  5.710 1.020 5.870 2.890 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.250 1.420 4.325 1.705 ;
        RECT  4.165 1.370 4.250 1.705 ;
        RECT  4.015 1.370 4.165 1.700 ;
        RECT  3.825 1.290 4.015 1.700 ;
        RECT  3.805 1.290 3.825 1.580 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 1.290 2.175 1.580 ;
        RECT  1.965 1.290 1.975 1.965 ;
        RECT  1.815 1.420 1.965 1.965 ;
        RECT  1.715 1.705 1.815 1.965 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.575 -0.250 6.900 0.250 ;
        RECT  6.315 -0.250 6.575 0.405 ;
        RECT  5.295 -0.250 6.315 0.250 ;
        RECT  5.035 -0.250 5.295 0.405 ;
        RECT  4.125 -0.250 5.035 0.250 ;
        RECT  3.865 -0.250 4.125 0.405 ;
        RECT  1.915 -0.250 3.865 0.250 ;
        RECT  1.655 -0.250 1.915 0.405 ;
        RECT  0.385 -0.250 1.655 0.250 ;
        RECT  0.125 -0.250 0.385 0.745 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.840 6.775 3.940 ;
        RECT  5.610 3.440 6.515 3.940 ;
        RECT  5.350 3.070 5.610 3.940 ;
        RECT  4.480 3.440 5.350 3.940 ;
        RECT  4.220 3.285 4.480 3.940 ;
        RECT  2.235 3.440 4.220 3.940 ;
        RECT  1.975 3.285 2.235 3.940 ;
        RECT  0.385 3.440 1.975 3.940 ;
        RECT  0.125 2.555 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.225 0.610 6.385 1.495 ;
        RECT  6.030 0.610 6.225 0.770 ;
        RECT  5.770 0.510 6.030 0.770 ;
        RECT  5.530 0.610 5.770 0.770 ;
        RECT  5.370 0.610 5.530 2.890 ;
        RECT  4.990 2.730 5.370 2.890 ;
        RECT  5.030 0.700 5.190 2.215 ;
        RECT  4.725 0.700 5.030 0.860 ;
        RECT  4.725 2.730 4.990 3.105 ;
        RECT  4.300 2.390 4.850 2.550 ;
        RECT  4.645 1.080 4.805 2.165 ;
        RECT  4.465 0.520 4.725 0.860 ;
        RECT  4.040 2.945 4.725 3.105 ;
        RECT  4.445 1.080 4.645 1.240 ;
        RECT  3.960 2.005 4.645 2.165 ;
        RECT  3.615 0.700 4.465 0.860 ;
        RECT  4.140 2.390 4.300 2.745 ;
        RECT  1.215 2.585 4.140 2.745 ;
        RECT  3.880 2.945 4.040 3.255 ;
        RECT  3.800 2.005 3.960 2.405 ;
        RECT  2.975 2.245 3.800 2.405 ;
        RECT  3.455 0.700 3.615 2.050 ;
        RECT  3.155 1.890 3.455 2.050 ;
        RECT  2.975 1.410 3.275 1.570 ;
        RECT  2.765 0.950 3.025 1.225 ;
        RECT  2.815 1.410 2.975 2.405 ;
        RECT  2.665 2.945 2.925 3.255 ;
        RECT  1.535 2.175 2.815 2.335 ;
        RECT  1.325 0.950 2.765 1.110 ;
        RECT  0.765 2.945 2.665 3.105 ;
        RECT  0.765 0.610 1.535 0.770 ;
        RECT  1.375 1.705 1.535 2.335 ;
        RECT  1.285 1.705 1.375 1.965 ;
        RECT  1.105 0.950 1.325 1.250 ;
        RECT  1.105 2.485 1.215 2.745 ;
        RECT  0.945 0.950 1.105 2.745 ;
        RECT  0.605 0.610 0.765 3.105 ;
        RECT  0.575 2.695 0.605 2.955 ;
    END
END TLATSRXL

MACRO TLATX4
    CLASS CORE ;
    FOREIGN TLATX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.025 1.700 7.235 2.400 ;
        RECT  6.795 1.700 7.025 2.395 ;
        RECT  6.775 1.055 6.795 2.395 ;
        RECT  6.725 1.055 6.775 2.585 ;
        RECT  6.555 0.695 6.725 3.010 ;
        RECT  6.465 0.695 6.555 1.295 ;
        RECT  6.465 2.070 6.555 3.010 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.705 1.290 5.855 2.220 ;
        RECT  5.445 0.695 5.705 2.220 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 0.880 0.370 1.895 ;
        RECT  0.110 1.515 0.125 1.895 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 1.485 1.835 1.990 ;
        RECT  1.505 1.700 1.575 1.990 ;
        END
        ANTENNAGATEAREA     0.4628 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 -0.250 7.360 0.250 ;
        RECT  6.975 -0.250 7.235 1.095 ;
        RECT  6.215 -0.250 6.975 0.250 ;
        RECT  5.955 -0.250 6.215 1.095 ;
        RECT  5.190 -0.250 5.955 0.250 ;
        RECT  4.930 -0.250 5.190 1.095 ;
        RECT  3.485 -0.250 4.930 0.250 ;
        RECT  3.225 -0.250 3.485 0.405 ;
        RECT  1.695 -0.250 3.225 0.250 ;
        RECT  1.435 -0.250 1.695 0.735 ;
        RECT  0.385 -0.250 1.435 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 3.440 7.360 3.940 ;
        RECT  6.975 2.600 7.235 3.940 ;
        RECT  6.215 3.440 6.975 3.940 ;
        RECT  5.955 2.940 6.215 3.940 ;
        RECT  5.165 3.440 5.955 3.940 ;
        RECT  4.905 3.285 5.165 3.940 ;
        RECT  3.415 3.440 4.905 3.940 ;
        RECT  3.155 3.285 3.415 3.940 ;
        RECT  1.580 3.440 3.155 3.940 ;
        RECT  1.320 2.955 1.580 3.940 ;
        RECT  0.385 3.440 1.320 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.260 1.580 6.360 1.840 ;
        RECT  6.100 1.580 6.260 2.760 ;
        RECT  5.225 2.600 6.100 2.760 ;
        RECT  5.065 1.275 5.225 2.760 ;
        RECT  4.750 1.275 5.065 1.440 ;
        RECT  4.705 2.600 5.065 2.760 ;
        RECT  4.405 1.620 4.885 1.780 ;
        RECT  4.610 0.655 4.750 1.440 ;
        RECT  4.545 2.250 4.705 2.940 ;
        RECT  4.590 0.550 4.610 1.440 ;
        RECT  4.350 0.550 4.590 0.815 ;
        RECT  3.270 2.780 4.545 2.940 ;
        RECT  4.365 1.110 4.405 2.050 ;
        RECT  4.245 1.110 4.365 2.600 ;
        RECT  3.985 0.655 4.350 0.815 ;
        RECT  2.585 1.110 4.245 1.270 ;
        RECT  4.205 1.890 4.245 2.600 ;
        RECT  2.560 2.440 4.205 2.600 ;
        RECT  3.940 1.480 4.065 1.640 ;
        RECT  3.725 0.470 3.985 0.815 ;
        RECT  3.780 1.480 3.940 2.260 ;
        RECT  2.315 2.100 3.780 2.260 ;
        RECT  2.795 1.760 3.585 1.920 ;
        RECT  2.635 1.465 2.795 1.920 ;
        RECT  2.535 1.465 2.635 1.745 ;
        RECT  2.375 0.685 2.585 1.285 ;
        RECT  2.435 2.440 2.560 2.775 ;
        RECT  2.175 1.465 2.535 1.625 ;
        RECT  2.400 2.440 2.435 3.215 ;
        RECT  2.175 2.615 2.400 3.215 ;
        RECT  2.325 0.685 2.375 0.945 ;
        RECT  2.215 1.805 2.315 2.260 ;
        RECT  2.055 1.805 2.215 2.335 ;
        RECT  2.015 1.140 2.175 1.625 ;
        RECT  1.605 2.175 2.055 2.335 ;
        RECT  1.265 1.140 2.015 1.300 ;
        RECT  1.445 2.175 1.605 2.775 ;
        RECT  0.785 2.615 1.445 2.775 ;
        RECT  1.255 1.140 1.265 2.400 ;
        RECT  1.105 0.525 1.255 2.400 ;
        RECT  1.095 0.525 1.105 1.300 ;
        RECT  0.925 2.140 1.105 2.400 ;
        RECT  0.925 0.525 1.095 0.785 ;
        RECT  0.710 1.640 0.925 1.900 ;
        RECT  0.710 1.035 0.815 1.295 ;
        RECT  0.710 2.615 0.785 2.910 ;
        RECT  0.550 1.035 0.710 2.910 ;
        RECT  0.525 2.650 0.550 2.910 ;
    END
END TLATX4

MACRO TLATX2
    CLASS CORE ;
    FOREIGN TLATX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 0.675 5.395 2.955 ;
        RECT  5.135 0.675 5.185 1.275 ;
        RECT  5.135 2.015 5.185 2.955 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.375 1.290 4.475 1.765 ;
        RECT  4.275 1.290 4.375 2.895 ;
        RECT  4.115 1.210 4.275 2.895 ;
        RECT  4.100 1.210 4.115 1.370 ;
        RECT  3.840 1.010 4.100 1.370 ;
        END
        ANTENNADIFFAREA     0.7458 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 0.880 0.370 1.975 ;
        RECT  0.110 1.715 0.125 1.975 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.395 1.865 1.655 ;
        RECT  1.715 1.395 1.765 1.985 ;
        RECT  1.605 1.395 1.715 1.990 ;
        RECT  1.505 1.700 1.605 1.990 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 -0.250 5.520 0.250 ;
        RECT  4.625 -0.250 4.885 0.685 ;
        RECT  3.395 -0.250 4.625 0.250 ;
        RECT  3.135 -0.250 3.395 0.405 ;
        RECT  1.605 -0.250 3.135 0.250 ;
        RECT  1.345 -0.250 1.605 0.405 ;
        RECT  0.385 -0.250 1.345 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 3.440 5.520 3.940 ;
        RECT  4.625 2.105 4.885 3.940 ;
        RECT  3.285 3.440 4.625 3.940 ;
        RECT  3.025 3.285 3.285 3.940 ;
        RECT  1.515 3.440 3.025 3.940 ;
        RECT  1.255 2.955 1.515 3.940 ;
        RECT  0.385 3.440 1.255 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.845 1.575 5.005 1.835 ;
        RECT  4.685 0.870 4.845 1.835 ;
        RECT  4.440 0.870 4.685 1.030 ;
        RECT  4.280 0.590 4.440 1.030 ;
        RECT  3.975 0.590 4.280 0.750 ;
        RECT  3.715 0.550 3.975 0.750 ;
        RECT  3.775 1.550 3.935 2.645 ;
        RECT  3.655 1.550 3.775 1.710 ;
        RECT  3.565 2.385 3.775 2.645 ;
        RECT  3.655 0.590 3.715 0.750 ;
        RECT  3.495 0.590 3.655 1.710 ;
        RECT  2.980 1.940 3.590 2.200 ;
        RECT  3.160 1.395 3.495 1.710 ;
        RECT  2.820 0.710 2.980 2.955 ;
        RECT  2.525 0.710 2.820 0.870 ;
        RECT  2.345 2.795 2.820 2.955 ;
        RECT  2.480 1.050 2.640 2.135 ;
        RECT  2.345 2.355 2.605 2.615 ;
        RECT  2.265 0.495 2.525 0.870 ;
        RECT  1.560 1.050 2.480 1.210 ;
        RECT  2.395 1.875 2.480 2.135 ;
        RECT  2.210 2.355 2.345 2.515 ;
        RECT  2.085 2.795 2.345 3.055 ;
        RECT  2.210 1.395 2.300 1.655 ;
        RECT  2.050 1.395 2.210 2.515 ;
        RECT  1.220 2.355 2.050 2.515 ;
        RECT  1.400 0.725 1.560 1.210 ;
        RECT  0.955 0.725 1.400 0.885 ;
        RECT  1.125 1.065 1.220 2.515 ;
        RECT  1.060 1.065 1.125 2.775 ;
        RECT  0.925 1.065 1.060 1.325 ;
        RECT  0.965 2.355 1.060 2.775 ;
        RECT  0.925 2.615 0.965 2.775 ;
        RECT  0.745 0.500 0.955 0.885 ;
        RECT  0.665 2.615 0.925 3.030 ;
        RECT  0.785 1.655 0.880 1.915 ;
        RECT  0.745 1.655 0.785 2.415 ;
        RECT  0.695 0.500 0.745 2.415 ;
        RECT  0.585 0.725 0.695 2.415 ;
        RECT  0.525 2.155 0.585 2.415 ;
    END
END TLATX2

MACRO TLATX1
    CLASS CORE ;
    FOREIGN TLATX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.425 1.515 4.475 2.585 ;
        RECT  4.415 1.515 4.425 2.715 ;
        RECT  4.265 1.025 4.415 2.715 ;
        RECT  4.255 1.025 4.265 2.335 ;
        END
        ANTENNADIFFAREA     0.4247 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.915 0.680 4.075 2.680 ;
        RECT  3.595 0.680 3.915 0.840 ;
        RECT  3.805 2.335 3.915 2.680 ;
        RECT  3.565 2.520 3.805 2.680 ;
        RECT  3.335 0.580 3.595 0.840 ;
        RECT  3.345 2.520 3.565 2.855 ;
        RECT  3.305 2.595 3.345 2.855 ;
        END
        ANTENNADIFFAREA     0.3796 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.475 0.445 1.735 ;
        RECT  0.125 1.120 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0676 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 1.700 1.715 1.990 ;
        RECT  1.505 1.180 1.555 1.990 ;
        RECT  1.395 1.180 1.505 1.925 ;
        END
        ANTENNAGATEAREA     0.1469 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 -0.250 4.600 0.250 ;
        RECT  3.940 -0.250 4.200 0.405 ;
        RECT  3.045 -0.250 3.940 0.250 ;
        RECT  2.785 -0.250 3.045 0.405 ;
        RECT  1.465 -0.250 2.785 0.250 ;
        RECT  1.205 -0.250 1.465 0.405 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 3.440 4.600 3.940 ;
        RECT  3.815 3.285 4.075 3.940 ;
        RECT  2.995 3.440 3.815 3.940 ;
        RECT  2.735 3.285 2.995 3.940 ;
        RECT  1.275 3.440 2.735 3.940 ;
        RECT  1.115 2.975 1.275 3.940 ;
        RECT  0.385 3.440 1.115 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.625 1.175 3.735 1.760 ;
        RECT  3.575 1.175 3.625 2.295 ;
        RECT  3.365 1.175 3.575 1.335 ;
        RECT  3.465 1.550 3.575 2.295 ;
        RECT  3.085 2.135 3.465 2.295 ;
        RECT  2.585 1.495 3.255 1.755 ;
        RECT  2.925 2.135 3.085 3.010 ;
        RECT  2.505 2.850 2.925 3.010 ;
        RECT  2.425 0.770 2.585 2.670 ;
        RECT  2.265 0.770 2.425 0.930 ;
        RECT  1.820 2.510 2.425 2.670 ;
        RECT  2.020 2.850 2.280 3.110 ;
        RECT  2.105 0.670 2.265 0.930 ;
        RECT  2.055 1.180 2.145 1.440 ;
        RECT  1.895 1.180 2.055 2.330 ;
        RECT  1.640 2.850 2.020 3.010 ;
        RECT  1.885 0.695 1.895 1.440 ;
        RECT  1.640 2.170 1.895 2.330 ;
        RECT  1.735 0.695 1.885 1.390 ;
        RECT  1.215 0.695 1.735 0.855 ;
        RECT  1.480 2.170 1.640 3.010 ;
        RECT  1.055 0.695 1.215 2.765 ;
        RECT  0.895 0.695 1.055 0.855 ;
        RECT  0.485 2.605 1.055 2.765 ;
        RECT  0.715 0.470 0.895 0.855 ;
        RECT  0.795 1.515 0.875 1.780 ;
        RECT  0.565 2.945 0.825 3.220 ;
        RECT  0.795 1.035 0.815 1.295 ;
        RECT  0.635 1.035 0.795 2.330 ;
        RECT  0.635 0.470 0.715 0.630 ;
        RECT  0.555 1.035 0.635 1.295 ;
        RECT  0.535 1.960 0.635 2.330 ;
        RECT  0.305 2.945 0.565 3.105 ;
        RECT  0.305 2.170 0.535 2.330 ;
        RECT  0.145 2.170 0.305 3.105 ;
    END
END TLATX1

MACRO TLATXL
    CLASS CORE ;
    FOREIGN TLATXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.425 1.515 4.475 2.810 ;
        RECT  4.265 1.025 4.425 2.810 ;
        RECT  4.205 2.305 4.265 2.810 ;
        END
        ANTENNADIFFAREA     0.2827 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.020 0.595 4.085 2.100 ;
        RECT  3.925 0.595 4.020 2.855 ;
        RECT  3.680 0.595 3.925 0.755 ;
        RECT  3.860 1.940 3.925 2.855 ;
        RECT  3.805 2.110 3.860 2.855 ;
        RECT  3.190 2.595 3.805 2.855 ;
        RECT  3.420 0.495 3.680 0.755 ;
        END
        ANTENNADIFFAREA     0.2340 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.475 0.445 1.735 ;
        RECT  0.125 1.120 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 1.700 1.715 1.990 ;
        RECT  1.505 1.120 1.555 1.990 ;
        RECT  1.395 1.120 1.505 1.925 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.280 -0.250 4.600 0.250 ;
        RECT  4.020 -0.250 4.280 0.405 ;
        RECT  3.095 -0.250 4.020 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  1.465 -0.250 2.835 0.250 ;
        RECT  1.205 -0.250 1.465 0.405 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.820 3.440 4.600 3.940 ;
        RECT  3.560 3.285 3.820 3.940 ;
        RECT  2.975 3.440 3.560 3.940 ;
        RECT  2.715 3.285 2.975 3.940 ;
        RECT  1.325 3.440 2.715 3.940 ;
        RECT  1.065 2.860 1.325 3.940 ;
        RECT  0.385 3.440 1.065 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.625 1.500 3.745 1.760 ;
        RECT  3.625 1.005 3.680 1.265 ;
        RECT  3.465 1.005 3.625 2.295 ;
        RECT  3.420 1.005 3.465 1.265 ;
        RECT  3.010 2.135 3.465 2.295 ;
        RECT  2.670 1.695 3.245 1.955 ;
        RECT  2.850 2.135 3.010 3.060 ;
        RECT  2.535 2.900 2.850 3.060 ;
        RECT  2.510 0.780 2.670 2.510 ;
        RECT  2.275 2.900 2.535 3.160 ;
        RECT  2.350 0.780 2.510 0.940 ;
        RECT  2.065 2.350 2.510 2.510 ;
        RECT  2.090 0.680 2.350 0.940 ;
        RECT  2.145 1.910 2.295 2.170 ;
        RECT  1.985 1.120 2.145 2.170 ;
        RECT  1.805 2.350 2.065 2.610 ;
        RECT  1.895 1.120 1.985 1.385 ;
        RECT  1.735 0.775 1.895 1.385 ;
        RECT  1.215 0.775 1.735 0.935 ;
        RECT  1.055 0.690 1.215 2.680 ;
        RECT  0.895 0.690 1.055 0.855 ;
        RECT  0.485 2.520 1.055 2.680 ;
        RECT  0.715 0.490 0.895 0.855 ;
        RECT  0.815 1.515 0.875 1.780 ;
        RECT  0.565 2.860 0.825 3.120 ;
        RECT  0.655 1.035 0.815 2.330 ;
        RECT  0.635 0.490 0.715 0.650 ;
        RECT  0.555 1.035 0.655 1.295 ;
        RECT  0.555 1.960 0.655 2.330 ;
        RECT  0.305 2.860 0.565 3.020 ;
        RECT  0.305 2.170 0.555 2.330 ;
        RECT  0.145 2.170 0.305 3.020 ;
    END
END TLATXL

MACRO SMDFFHQX8
    CLASS CORE ;
    FOREIGN SMDFFHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.540 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.105 1.335 6.615 1.495 ;
        RECT  5.945 0.585 6.105 1.495 ;
        RECT  3.790 0.585 5.945 0.745 ;
        RECT  3.630 0.470 3.790 0.745 ;
        RECT  1.530 0.470 3.630 0.630 ;
        RECT  1.525 0.470 1.530 0.695 ;
        RECT  1.245 0.430 1.525 0.745 ;
        RECT  1.230 0.535 1.245 0.745 ;
        RECT  0.795 0.585 1.230 0.745 ;
        RECT  0.715 0.585 0.795 1.680 ;
        RECT  0.635 0.585 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.745 7.185 1.905 ;
        RECT  5.850 1.700 5.855 1.990 ;
        RECT  5.645 1.675 5.850 1.990 ;
        RECT  5.485 1.575 5.645 1.835 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.900 1.105 21.955 2.585 ;
        RECT  21.640 0.695 21.900 2.895 ;
        RECT  21.035 1.290 21.640 1.990 ;
        RECT  20.875 1.290 21.035 2.175 ;
        RECT  20.615 0.695 20.875 2.895 ;
        END
        ANTENNADIFFAREA     1.5960 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.670 2.805 2.030 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.325 1.185 9.640 1.680 ;
        END
        ANTENNAGATEAREA     0.2730 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  10.915 1.160 11.360 1.420 ;
        RECT  10.705 1.160 10.915 1.580 ;
        RECT  10.420 1.160 10.705 1.420 ;
        END
        ANTENNAGATEAREA     0.4238 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.410 -0.250 22.540 0.250 ;
        RECT  22.150 -0.250 22.410 1.115 ;
        RECT  21.385 -0.250 22.150 0.250 ;
        RECT  21.125 -0.250 21.385 1.065 ;
        RECT  20.325 -0.250 21.125 0.250 ;
        RECT  20.065 -0.250 20.325 0.405 ;
        RECT  19.445 -0.250 20.065 0.250 ;
        RECT  19.185 -0.250 19.445 0.405 ;
        RECT  16.610 -0.250 19.185 0.250 ;
        RECT  16.350 -0.250 16.610 0.785 ;
        RECT  15.530 -0.250 16.350 0.250 ;
        RECT  15.270 -0.250 15.530 0.865 ;
        RECT  14.420 -0.250 15.270 0.250 ;
        RECT  14.160 -0.250 14.420 0.405 ;
        RECT  12.690 -0.250 14.160 0.250 ;
        RECT  12.430 -0.250 12.690 0.405 ;
        RECT  11.405 -0.250 12.430 0.250 ;
        RECT  11.145 -0.250 11.405 0.405 ;
        RECT  10.325 -0.250 11.145 0.250 ;
        RECT  10.065 -0.250 10.325 0.405 ;
        RECT  9.275 -0.250 10.065 0.250 ;
        RECT  9.015 -0.250 9.275 0.405 ;
        RECT  7.375 -0.250 9.015 0.250 ;
        RECT  7.115 -0.250 7.375 0.405 ;
        RECT  6.235 -0.250 7.115 0.250 ;
        RECT  5.975 -0.250 6.235 0.405 ;
        RECT  4.235 -0.250 5.975 0.250 ;
        RECT  3.975 -0.250 4.235 0.405 ;
        RECT  0.815 -0.250 3.975 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.410 3.440 22.540 3.940 ;
        RECT  22.150 2.255 22.410 3.940 ;
        RECT  21.385 3.440 22.150 3.940 ;
        RECT  21.125 2.595 21.385 3.940 ;
        RECT  20.360 3.440 21.125 3.940 ;
        RECT  20.100 2.935 20.360 3.940 ;
        RECT  19.455 3.440 20.100 3.940 ;
        RECT  19.195 2.475 19.455 3.940 ;
        RECT  16.895 3.440 19.195 3.940 ;
        RECT  16.635 3.285 16.895 3.940 ;
        RECT  15.815 3.440 16.635 3.940 ;
        RECT  15.555 3.285 15.815 3.940 ;
        RECT  14.545 3.440 15.555 3.940 ;
        RECT  14.285 2.890 14.545 3.940 ;
        RECT  12.835 3.440 14.285 3.940 ;
        RECT  12.575 3.285 12.835 3.940 ;
        RECT  11.745 3.440 12.575 3.940 ;
        RECT  11.485 3.285 11.745 3.940 ;
        RECT  9.795 3.440 11.485 3.940 ;
        RECT  9.535 3.285 9.795 3.940 ;
        RECT  7.695 3.440 9.535 3.940 ;
        RECT  7.435 3.285 7.695 3.940 ;
        RECT  6.645 3.440 7.435 3.940 ;
        RECT  6.385 2.945 6.645 3.940 ;
        RECT  5.490 3.440 6.385 3.940 ;
        RECT  5.230 3.285 5.490 3.940 ;
        RECT  4.285 3.405 5.230 3.940 ;
        RECT  4.025 3.095 4.285 3.940 ;
        RECT  0.815 3.440 4.025 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.330 1.490 20.430 1.750 ;
        RECT  20.170 0.605 20.330 1.750 ;
        RECT  18.540 0.605 20.170 0.765 ;
        RECT  19.915 2.425 19.965 2.685 ;
        RECT  19.755 0.945 19.915 2.685 ;
        RECT  19.650 0.945 19.755 1.105 ;
        RECT  19.185 1.555 19.755 1.845 ;
        RECT  19.705 2.425 19.755 2.685 ;
        RECT  18.845 1.055 19.005 3.100 ;
        RECT  18.710 1.055 18.845 1.215 ;
        RECT  14.985 2.940 18.845 3.100 ;
        RECT  18.550 0.955 18.710 1.215 ;
        RECT  18.505 1.955 18.665 2.215 ;
        RECT  18.370 0.515 18.540 0.775 ;
        RECT  18.370 1.955 18.505 2.115 ;
        RECT  18.210 0.515 18.370 2.115 ;
        RECT  18.055 2.465 18.315 2.725 ;
        RECT  17.520 0.665 18.210 0.830 ;
        RECT  17.805 1.955 18.210 2.115 ;
        RECT  17.295 2.565 18.055 2.725 ;
        RECT  17.930 1.035 18.030 1.295 ;
        RECT  17.770 1.035 17.930 1.605 ;
        RECT  17.545 1.955 17.805 2.215 ;
        RECT  17.245 1.445 17.770 1.605 ;
        RECT  17.260 0.665 17.520 1.265 ;
        RECT  17.245 2.125 17.295 2.725 ;
        RECT  17.085 1.445 17.245 2.725 ;
        RECT  17.015 1.445 17.085 1.605 ;
        RECT  17.035 2.125 17.085 2.725 ;
        RECT  16.355 2.565 17.035 2.725 ;
        RECT  16.855 1.035 17.015 1.605 ;
        RECT  16.750 1.035 16.855 1.295 ;
        RECT  16.070 1.135 16.750 1.295 ;
        RECT  15.320 1.585 16.525 1.845 ;
        RECT  16.095 2.125 16.355 2.725 ;
        RECT  15.585 2.360 16.095 2.520 ;
        RECT  15.810 0.690 16.070 1.295 ;
        RECT  15.325 2.360 15.585 2.620 ;
        RECT  15.160 1.135 15.320 2.180 ;
        RECT  14.790 1.135 15.160 1.295 ;
        RECT  14.905 2.020 15.160 2.180 ;
        RECT  14.730 0.535 14.990 0.795 ;
        RECT  14.825 2.550 14.985 3.100 ;
        RECT  14.645 2.020 14.905 2.280 ;
        RECT  14.090 2.550 14.825 2.710 ;
        RECT  14.530 1.035 14.790 1.295 ;
        RECT  13.935 0.585 14.730 0.745 ;
        RECT  14.420 1.475 14.680 1.735 ;
        RECT  13.685 2.020 14.645 2.180 ;
        RECT  13.585 1.085 14.530 1.245 ;
        RECT  13.245 1.475 14.420 1.635 ;
        RECT  13.930 2.550 14.090 2.765 ;
        RECT  13.775 0.480 13.935 0.745 ;
        RECT  13.245 2.605 13.930 2.765 ;
        RECT  13.255 2.945 13.855 3.215 ;
        RECT  13.060 0.480 13.775 0.640 ;
        RECT  13.425 2.020 13.685 2.280 ;
        RECT  13.425 0.820 13.585 1.245 ;
        RECT  13.310 0.820 13.425 0.980 ;
        RECT  8.695 2.945 13.255 3.105 ;
        RECT  13.085 1.245 13.245 2.765 ;
        RECT  12.920 1.245 13.085 1.405 ;
        RECT  9.980 2.605 13.085 2.765 ;
        RECT  12.900 0.480 13.060 0.920 ;
        RECT  12.660 1.145 12.920 1.405 ;
        RECT  12.470 1.610 12.905 1.885 ;
        RECT  12.470 0.760 12.900 0.920 ;
        RECT  12.310 0.760 12.470 2.285 ;
        RECT  11.890 0.885 12.310 1.145 ;
        RECT  12.295 2.125 12.310 2.285 ;
        RECT  12.035 2.125 12.295 2.385 ;
        RECT  11.700 1.650 12.125 1.935 ;
        RECT  10.335 2.225 12.035 2.385 ;
        RECT  11.540 0.710 11.700 1.935 ;
        RECT  10.865 0.710 11.540 0.870 ;
        RECT  10.545 1.775 11.540 1.935 ;
        RECT  10.605 0.610 10.865 0.870 ;
        RECT  10.285 1.775 10.545 2.040 ;
        RECT  9.820 0.710 9.980 2.765 ;
        RECT  9.785 0.710 9.820 0.870 ;
        RECT  9.525 0.610 9.785 0.870 ;
        RECT  9.140 1.955 9.255 2.555 ;
        RECT  8.995 0.745 9.140 2.555 ;
        RECT  8.980 0.745 8.995 2.120 ;
        RECT  8.735 0.745 8.980 0.905 ;
        RECT  8.475 0.645 8.735 0.905 ;
        RECT  8.535 1.085 8.695 3.105 ;
        RECT  8.295 1.085 8.535 1.245 ;
        RECT  7.135 2.945 8.535 3.105 ;
        RECT  8.265 1.425 8.325 2.715 ;
        RECT  8.225 0.595 8.295 1.245 ;
        RECT  8.165 1.425 8.265 2.765 ;
        RECT  8.135 0.495 8.225 1.245 ;
        RECT  7.955 1.425 8.165 1.585 ;
        RECT  8.005 2.505 8.165 2.765 ;
        RECT  7.965 0.495 8.135 0.755 ;
        RECT  7.795 1.055 7.955 1.585 ;
        RECT  7.615 1.795 7.895 2.055 ;
        RECT  7.565 1.055 7.795 1.215 ;
        RECT  7.455 1.395 7.615 2.275 ;
        RECT  7.385 1.395 7.455 1.555 ;
        RECT  7.095 2.115 7.455 2.275 ;
        RECT  7.225 0.995 7.385 1.555 ;
        RECT  6.815 0.995 7.225 1.155 ;
        RECT  6.975 2.520 7.135 3.105 ;
        RECT  4.965 2.520 6.975 2.680 ;
        RECT  6.555 0.895 6.815 1.155 ;
        RECT  4.625 2.860 6.185 3.020 ;
        RECT  5.305 2.170 6.065 2.330 ;
        RECT  5.305 1.045 5.495 1.305 ;
        RECT  5.235 1.045 5.305 2.330 ;
        RECT  5.145 1.145 5.235 2.330 ;
        RECT  4.575 1.635 5.145 1.895 ;
        RECT  4.805 2.415 4.965 2.680 ;
        RECT  4.395 0.925 4.815 1.085 ;
        RECT  4.055 2.415 4.805 2.575 ;
        RECT  4.395 2.075 4.760 2.235 ;
        RECT  4.465 2.755 4.625 3.020 ;
        RECT  3.825 2.755 4.465 2.915 ;
        RECT  4.235 0.925 4.395 2.235 ;
        RECT  3.435 0.925 4.235 1.085 ;
        RECT  3.895 1.400 4.055 2.575 ;
        RECT  3.840 1.400 3.895 1.560 ;
        RECT  3.485 2.415 3.895 2.575 ;
        RECT  3.580 1.300 3.840 1.560 ;
        RECT  3.665 2.755 3.825 3.220 ;
        RECT  1.200 3.060 3.665 3.220 ;
        RECT  3.325 2.415 3.485 2.880 ;
        RECT  3.275 0.810 3.435 1.085 ;
        RECT  1.710 2.720 3.325 2.880 ;
        RECT  3.145 1.300 3.315 1.560 ;
        RECT  2.065 0.925 3.275 1.085 ;
        RECT  3.055 1.300 3.145 2.480 ;
        RECT  2.985 1.350 3.055 2.480 ;
        RECT  2.245 2.220 2.985 2.380 ;
        RECT  2.195 1.320 2.275 1.480 ;
        RECT  2.195 2.220 2.245 2.480 ;
        RECT  2.035 1.320 2.195 2.480 ;
        RECT  1.905 0.810 2.065 1.085 ;
        RECT  2.015 1.320 2.035 1.480 ;
        RECT  1.985 2.220 2.035 2.480 ;
        RECT  1.710 1.210 1.760 1.470 ;
        RECT  1.550 1.210 1.710 2.880 ;
        RECT  1.500 1.210 1.550 1.470 ;
        RECT  1.445 2.420 1.550 2.680 ;
        RECT  1.040 2.580 1.200 3.220 ;
        RECT  0.385 2.580 1.040 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.125 1.025 0.225 2.515 ;
        RECT  0.115 1.035 0.125 2.515 ;
    END
END SMDFFHQX8

MACRO SMDFFHQX4
    CLASS CORE ;
    FOREIGN SMDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.160 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.105 1.345 6.445 1.505 ;
        RECT  5.945 0.585 6.105 1.505 ;
        RECT  3.760 0.585 5.945 0.745 ;
        RECT  3.600 0.470 3.760 0.745 ;
        RECT  1.530 0.470 3.600 0.630 ;
        RECT  1.525 0.470 1.530 0.695 ;
        RECT  1.245 0.430 1.525 0.745 ;
        RECT  1.230 0.535 1.245 0.745 ;
        RECT  0.795 0.585 1.230 0.745 ;
        RECT  0.635 0.585 0.795 1.580 ;
        RECT  0.585 1.105 0.635 1.580 ;
        RECT  0.455 1.315 0.585 1.575 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 1.745 7.015 1.905 ;
        RECT  6.105 1.700 6.315 1.990 ;
        RECT  5.485 1.700 6.105 1.870 ;
        RECT  5.325 1.575 5.485 1.870 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.525 1.105 20.575 2.585 ;
        RECT  20.515 0.695 20.525 2.585 ;
        RECT  20.265 0.695 20.515 2.895 ;
        RECT  20.255 1.510 20.265 2.895 ;
        END
        ANTENNADIFFAREA     0.7980 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.670 2.805 2.030 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.325 1.290 9.535 1.670 ;
        RECT  9.045 1.335 9.325 1.670 ;
        END
        ANTENNAGATEAREA     0.2730 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  10.455 1.160 10.680 1.420 ;
        RECT  10.245 1.160 10.455 1.580 ;
        RECT  10.080 1.160 10.245 1.420 ;
        END
        ANTENNAGATEAREA     0.4238 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.035 -0.250 21.160 0.250 ;
        RECT  20.775 -0.250 21.035 1.115 ;
        RECT  19.975 -0.250 20.775 0.250 ;
        RECT  19.715 -0.250 19.975 0.405 ;
        RECT  19.175 -0.250 19.715 0.250 ;
        RECT  18.915 -0.250 19.175 0.405 ;
        RECT  16.385 -0.250 18.915 0.250 ;
        RECT  16.125 -0.250 16.385 0.785 ;
        RECT  15.275 -0.250 16.125 0.250 ;
        RECT  15.015 -0.250 15.275 0.865 ;
        RECT  14.000 -0.250 15.015 0.250 ;
        RECT  13.740 -0.250 14.000 0.405 ;
        RECT  12.255 -0.250 13.740 0.250 ;
        RECT  11.995 -0.250 12.255 0.405 ;
        RECT  11.310 -0.250 11.995 0.250 ;
        RECT  11.050 -0.250 11.310 0.405 ;
        RECT  10.230 -0.250 11.050 0.250 ;
        RECT  9.970 -0.250 10.230 0.405 ;
        RECT  9.020 -0.250 9.970 0.250 ;
        RECT  8.760 -0.250 9.020 0.405 ;
        RECT  7.140 -0.250 8.760 0.250 ;
        RECT  6.880 -0.250 7.140 0.405 ;
        RECT  6.075 -0.250 6.880 0.250 ;
        RECT  5.815 -0.250 6.075 0.405 ;
        RECT  4.200 -0.250 5.815 0.250 ;
        RECT  3.940 -0.250 4.200 0.405 ;
        RECT  0.815 -0.250 3.940 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.025 3.440 21.160 3.940 ;
        RECT  20.765 2.255 21.025 3.940 ;
        RECT  20.005 3.440 20.765 3.940 ;
        RECT  19.745 2.935 20.005 3.940 ;
        RECT  19.095 3.440 19.745 3.940 ;
        RECT  18.835 2.385 19.095 3.940 ;
        RECT  16.535 3.440 18.835 3.940 ;
        RECT  16.275 3.285 16.535 3.940 ;
        RECT  14.345 3.440 16.275 3.940 ;
        RECT  14.085 3.285 14.345 3.940 ;
        RECT  12.645 3.440 14.085 3.940 ;
        RECT  12.385 3.285 12.645 3.940 ;
        RECT  11.565 3.440 12.385 3.940 ;
        RECT  11.305 3.285 11.565 3.940 ;
        RECT  9.625 3.440 11.305 3.940 ;
        RECT  9.365 3.285 9.625 3.940 ;
        RECT  7.345 3.440 9.365 3.940 ;
        RECT  7.085 3.285 7.345 3.940 ;
        RECT  6.475 3.440 7.085 3.940 ;
        RECT  6.215 2.945 6.475 3.940 ;
        RECT  5.330 3.440 6.215 3.940 ;
        RECT  5.070 3.285 5.330 3.940 ;
        RECT  4.285 3.405 5.070 3.940 ;
        RECT  4.025 3.095 4.285 3.940 ;
        RECT  0.815 3.440 4.025 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.010 1.490 20.055 1.750 ;
        RECT  19.850 0.585 20.010 1.750 ;
        RECT  18.235 0.585 19.850 0.745 ;
        RECT  19.795 1.490 19.850 1.750 ;
        RECT  19.555 0.925 19.605 1.085 ;
        RECT  19.555 2.390 19.605 2.650 ;
        RECT  19.395 0.925 19.555 2.650 ;
        RECT  19.345 0.925 19.395 1.085 ;
        RECT  18.985 1.555 19.395 1.715 ;
        RECT  19.345 2.390 19.395 2.650 ;
        RECT  18.825 1.555 18.985 1.820 ;
        RECT  18.485 1.035 18.645 3.100 ;
        RECT  18.435 1.035 18.485 1.195 ;
        RECT  15.585 2.940 18.485 3.100 ;
        RECT  18.275 0.930 18.435 1.195 ;
        RECT  18.145 1.955 18.305 2.215 ;
        RECT  18.095 0.485 18.235 0.745 ;
        RECT  18.095 1.955 18.145 2.115 ;
        RECT  17.975 0.485 18.095 2.115 ;
        RECT  17.935 0.585 17.975 2.115 ;
        RECT  17.695 2.465 17.955 2.725 ;
        RECT  17.295 0.585 17.935 0.745 ;
        RECT  17.445 1.955 17.935 2.115 ;
        RECT  17.595 1.035 17.755 1.605 ;
        RECT  16.935 2.565 17.695 2.725 ;
        RECT  16.835 1.445 17.595 1.605 ;
        RECT  17.185 1.955 17.445 2.215 ;
        RECT  17.035 0.585 17.295 1.265 ;
        RECT  16.835 2.125 16.935 2.725 ;
        RECT  16.675 1.035 16.835 2.725 ;
        RECT  15.845 1.035 16.675 1.295 ;
        RECT  15.995 2.565 16.675 2.725 ;
        RECT  14.940 1.585 16.120 1.845 ;
        RECT  15.735 2.125 15.995 2.725 ;
        RECT  15.585 0.690 15.845 1.295 ;
        RECT  15.155 2.565 15.735 2.725 ;
        RECT  15.425 2.940 15.585 3.190 ;
        RECT  14.715 3.030 15.425 3.190 ;
        RECT  14.945 2.565 15.155 2.850 ;
        RECT  14.895 2.690 14.945 2.850 ;
        RECT  14.780 1.135 14.940 2.180 ;
        RECT  14.565 1.135 14.780 1.295 ;
        RECT  14.665 2.020 14.780 2.180 ;
        RECT  14.505 0.535 14.765 0.795 ;
        RECT  14.665 2.605 14.715 2.765 ;
        RECT  14.555 2.945 14.715 3.190 ;
        RECT  14.505 2.020 14.665 2.765 ;
        RECT  14.305 1.035 14.565 1.295 ;
        RECT  14.005 2.945 14.555 3.105 ;
        RECT  13.475 0.585 14.505 0.745 ;
        RECT  13.495 2.020 14.505 2.180 ;
        RECT  14.455 2.605 14.505 2.765 ;
        RECT  14.195 1.475 14.455 1.735 ;
        RECT  14.265 1.035 14.305 1.195 ;
        RECT  14.105 0.925 14.265 1.195 ;
        RECT  13.045 1.475 14.195 1.635 ;
        RECT  13.135 0.925 14.105 1.085 ;
        RECT  13.845 2.605 14.005 3.105 ;
        RECT  13.045 2.605 13.845 2.765 ;
        RECT  13.065 2.945 13.665 3.215 ;
        RECT  13.235 2.020 13.495 2.280 ;
        RECT  13.315 0.485 13.475 0.745 ;
        RECT  12.595 0.485 13.315 0.645 ;
        RECT  12.875 0.825 13.135 1.085 ;
        RECT  8.525 2.945 13.065 3.105 ;
        RECT  12.885 1.285 13.045 2.765 ;
        RECT  12.435 1.285 12.885 1.445 ;
        RECT  9.875 2.605 12.885 2.765 ;
        RECT  12.105 1.625 12.705 1.885 ;
        RECT  12.435 0.485 12.595 0.745 ;
        RECT  12.095 0.585 12.435 0.745 ;
        RECT  12.275 1.145 12.435 1.445 ;
        RECT  12.095 1.625 12.105 2.385 ;
        RECT  11.935 0.585 12.095 2.385 ;
        RECT  11.455 0.885 11.935 1.145 ;
        RECT  11.845 2.125 11.935 2.385 ;
        RECT  10.165 2.225 11.845 2.385 ;
        RECT  11.080 1.650 11.755 1.935 ;
        RECT  10.920 0.710 11.080 1.935 ;
        RECT  10.770 0.710 10.920 0.870 ;
        RECT  10.215 1.775 10.920 1.935 ;
        RECT  10.510 0.610 10.770 0.870 ;
        RECT  10.055 1.775 10.215 2.040 ;
        RECT  9.715 0.710 9.875 2.765 ;
        RECT  9.690 0.710 9.715 0.870 ;
        RECT  9.430 0.610 9.690 0.870 ;
        RECT  8.865 1.955 9.085 2.555 ;
        RECT  8.825 0.675 8.865 2.555 ;
        RECT  8.705 0.675 8.825 2.120 ;
        RECT  8.480 0.675 8.705 0.835 ;
        RECT  8.365 1.015 8.525 3.105 ;
        RECT  8.220 0.575 8.480 0.835 ;
        RECT  8.040 1.015 8.365 1.175 ;
        RECT  6.830 2.945 8.365 3.105 ;
        RECT  7.970 0.595 8.040 1.175 ;
        RECT  7.880 0.495 7.970 1.175 ;
        RECT  7.765 1.360 7.925 2.765 ;
        RECT  7.710 0.495 7.880 0.755 ;
        RECT  7.695 1.360 7.765 1.520 ;
        RECT  7.665 2.505 7.765 2.765 ;
        RECT  7.535 1.055 7.695 1.520 ;
        RECT  7.310 1.055 7.535 1.215 ;
        RECT  7.355 1.695 7.445 2.055 ;
        RECT  7.195 1.400 7.355 2.275 ;
        RECT  6.800 1.400 7.195 1.560 ;
        RECT  6.925 2.115 7.195 2.275 ;
        RECT  6.670 2.520 6.830 3.105 ;
        RECT  6.640 0.995 6.800 1.560 ;
        RECT  4.965 2.520 6.670 2.680 ;
        RECT  6.535 0.995 6.640 1.155 ;
        RECT  6.535 0.490 6.585 0.750 ;
        RECT  6.375 0.490 6.535 1.155 ;
        RECT  6.325 0.490 6.375 0.750 ;
        RECT  4.625 2.860 6.030 3.020 ;
        RECT  5.800 2.170 5.905 2.330 ;
        RECT  5.640 2.055 5.800 2.330 ;
        RECT  5.140 2.055 5.640 2.215 ;
        RECT  5.140 1.045 5.335 1.305 ;
        RECT  5.075 1.045 5.140 2.215 ;
        RECT  4.980 1.145 5.075 2.215 ;
        RECT  4.415 1.635 4.980 1.895 ;
        RECT  4.805 2.415 4.965 2.680 ;
        RECT  3.740 2.415 4.805 2.575 ;
        RECT  4.225 0.925 4.780 1.085 ;
        RECT  4.225 2.075 4.760 2.235 ;
        RECT  4.465 2.755 4.625 3.020 ;
        RECT  3.825 2.755 4.465 2.915 ;
        RECT  4.065 0.925 4.225 2.235 ;
        RECT  3.420 0.925 4.065 1.085 ;
        RECT  3.740 1.300 3.840 1.560 ;
        RECT  3.665 2.755 3.825 3.220 ;
        RECT  3.580 1.300 3.740 2.575 ;
        RECT  1.200 3.060 3.665 3.220 ;
        RECT  3.485 2.415 3.580 2.575 ;
        RECT  3.325 2.415 3.485 2.880 ;
        RECT  3.260 0.810 3.420 1.085 ;
        RECT  1.710 2.720 3.325 2.880 ;
        RECT  3.145 1.300 3.315 1.560 ;
        RECT  2.065 0.925 3.260 1.085 ;
        RECT  3.055 1.300 3.145 2.480 ;
        RECT  2.985 1.350 3.055 2.480 ;
        RECT  2.245 2.220 2.985 2.380 ;
        RECT  2.175 1.320 2.275 1.480 ;
        RECT  2.175 2.220 2.245 2.480 ;
        RECT  2.015 1.320 2.175 2.480 ;
        RECT  1.905 0.810 2.065 1.085 ;
        RECT  1.985 2.220 2.015 2.480 ;
        RECT  1.710 1.210 1.760 1.470 ;
        RECT  1.550 1.210 1.710 2.880 ;
        RECT  1.500 1.210 1.550 1.470 ;
        RECT  1.445 2.420 1.550 2.680 ;
        RECT  1.040 2.580 1.200 3.220 ;
        RECT  0.385 2.580 1.040 2.740 ;
        RECT  0.275 0.875 0.385 1.135 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 0.875 0.275 2.740 ;
        RECT  0.115 0.875 0.225 2.515 ;
    END
END SMDFFHQX4

MACRO SMDFFHQX2
    CLASS CORE ;
    FOREIGN SMDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.640 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.115 1.335 5.450 1.495 ;
        RECT  4.955 0.935 5.115 1.495 ;
        RECT  4.520 0.935 4.955 1.095 ;
        RECT  4.360 0.620 4.520 1.095 ;
        RECT  2.955 0.620 4.360 0.780 ;
        RECT  2.795 0.490 2.955 0.780 ;
        RECT  2.500 0.490 2.795 0.650 ;
        RECT  2.340 0.430 2.500 0.650 ;
        RECT  1.675 0.430 2.340 0.590 ;
        RECT  1.515 0.430 1.675 0.785 ;
        RECT  0.795 0.625 1.515 0.785 ;
        RECT  0.715 0.625 0.795 1.680 ;
        RECT  0.635 0.625 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 1.725 5.930 1.885 ;
        RECT  4.930 1.700 4.935 1.990 ;
        RECT  4.725 1.675 4.930 1.990 ;
        RECT  4.285 1.675 4.725 1.835 ;
        RECT  4.125 1.575 4.285 1.835 ;
        END
        ANTENNAGATEAREA     0.1001 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.255 0.695 15.515 2.895 ;
        END
        ANTENNADIFFAREA     0.7140 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.535 2.635 1.990 ;
        RECT  2.305 1.535 2.425 1.895 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.260 1.290 8.615 1.580 ;
        RECT  8.000 1.290 8.260 1.610 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.530 1.290 9.535 1.580 ;
        RECT  9.135 1.290 9.530 1.600 ;
        END
        ANTENNAGATEAREA     0.2327 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.975 -0.250 15.640 0.250 ;
        RECT  14.715 -0.250 14.975 0.405 ;
        RECT  14.175 -0.250 14.715 0.250 ;
        RECT  13.915 -0.250 14.175 0.405 ;
        RECT  12.055 -0.250 13.915 0.250 ;
        RECT  11.795 -0.250 12.055 0.755 ;
        RECT  10.405 -0.250 11.795 0.250 ;
        RECT  10.145 -0.250 10.405 0.405 ;
        RECT  8.800 -0.250 10.145 0.250 ;
        RECT  7.780 -0.250 8.800 0.405 ;
        RECT  6.140 -0.250 7.780 0.250 ;
        RECT  5.880 -0.250 6.140 0.405 ;
        RECT  4.990 -0.250 5.880 0.250 ;
        RECT  4.730 -0.250 4.990 0.745 ;
        RECT  3.395 -0.250 4.730 0.250 ;
        RECT  3.135 -0.250 3.395 0.405 ;
        RECT  0.815 -0.250 3.135 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.975 3.440 15.640 3.940 ;
        RECT  14.715 2.890 14.975 3.940 ;
        RECT  14.125 3.440 14.715 3.940 ;
        RECT  13.865 2.890 14.125 3.940 ;
        RECT  12.195 3.440 13.865 3.940 ;
        RECT  11.935 3.285 12.195 3.940 ;
        RECT  10.435 3.440 11.935 3.940 ;
        RECT  10.175 3.285 10.435 3.940 ;
        RECT  8.415 3.440 10.175 3.940 ;
        RECT  8.155 3.285 8.415 3.940 ;
        RECT  6.485 3.440 8.155 3.940 ;
        RECT  6.225 3.285 6.485 3.940 ;
        RECT  5.250 3.440 6.225 3.940 ;
        RECT  4.990 2.925 5.250 3.940 ;
        RECT  4.165 3.440 4.990 3.940 ;
        RECT  3.905 3.285 4.165 3.940 ;
        RECT  3.235 3.440 3.905 3.940 ;
        RECT  3.075 3.035 3.235 3.940 ;
        RECT  0.815 3.440 3.075 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.555 2.105 14.605 2.365 ;
        RECT  14.395 1.035 14.555 2.365 ;
        RECT  14.345 2.005 14.395 2.365 ;
        RECT  13.875 2.005 14.345 2.165 ;
        RECT  14.055 0.585 14.215 1.665 ;
        RECT  13.105 0.585 14.055 0.745 ;
        RECT  13.715 1.885 13.875 2.165 ;
        RECT  13.535 2.920 13.615 3.180 ;
        RECT  13.375 0.925 13.535 3.180 ;
        RECT  13.265 0.925 13.375 1.190 ;
        RECT  13.355 2.860 13.375 3.180 ;
        RECT  11.510 2.860 13.355 3.020 ;
        RECT  13.085 1.440 13.195 2.555 ;
        RECT  13.085 0.535 13.105 0.795 ;
        RECT  13.035 0.535 13.085 2.555 ;
        RECT  12.925 0.535 13.035 1.600 ;
        RECT  12.845 0.535 12.925 0.795 ;
        RECT  12.595 1.085 12.735 2.675 ;
        RECT  12.575 0.985 12.595 2.675 ;
        RECT  12.335 0.985 12.575 1.245 ;
        RECT  12.475 2.075 12.575 2.675 ;
        RECT  11.965 2.515 12.475 2.675 ;
        RECT  12.120 1.585 12.345 1.845 ;
        RECT  11.960 1.025 12.120 2.230 ;
        RECT  11.705 2.415 11.965 2.675 ;
        RECT  11.315 1.025 11.960 1.185 ;
        RECT  11.025 2.070 11.960 2.230 ;
        RECT  10.215 0.585 11.515 0.745 ;
        RECT  11.350 2.605 11.510 3.020 ;
        RECT  10.845 1.615 11.485 1.875 ;
        RECT  10.845 2.605 11.350 2.765 ;
        RECT  11.055 0.925 11.315 1.185 ;
        RECT  11.020 3.100 11.115 3.260 ;
        RECT  10.855 2.945 11.020 3.260 ;
        RECT  7.435 2.945 10.855 3.105 ;
        RECT  10.685 1.270 10.845 2.765 ;
        RECT  10.555 1.270 10.685 1.430 ;
        RECT  8.775 2.605 10.685 2.765 ;
        RECT  10.395 1.170 10.555 1.430 ;
        RECT  10.215 1.650 10.505 1.910 ;
        RECT  10.055 0.585 10.215 2.385 ;
        RECT  9.865 0.585 10.055 0.770 ;
        RECT  8.955 2.225 10.055 2.385 ;
        RECT  9.715 0.950 9.875 1.940 ;
        RECT  9.605 0.510 9.865 0.770 ;
        RECT  9.300 0.950 9.715 1.110 ;
        RECT  9.295 1.780 9.715 1.940 ;
        RECT  9.140 0.840 9.300 1.110 ;
        RECT  9.135 1.780 9.295 2.040 ;
        RECT  8.795 0.940 8.955 1.920 ;
        RECT  8.400 0.940 8.795 1.100 ;
        RECT  8.775 1.760 8.795 1.920 ;
        RECT  8.615 1.760 8.775 2.765 ;
        RECT  8.140 0.840 8.400 1.100 ;
        RECT  7.775 1.955 7.995 2.555 ;
        RECT  7.735 0.670 7.775 2.555 ;
        RECT  7.615 0.670 7.735 2.120 ;
        RECT  7.230 0.670 7.615 0.830 ;
        RECT  7.275 1.085 7.435 3.105 ;
        RECT  7.050 1.085 7.275 1.245 ;
        RECT  6.095 2.945 7.275 3.105 ;
        RECT  6.905 1.425 7.065 2.765 ;
        RECT  6.890 0.455 7.050 1.245 ;
        RECT  6.710 1.425 6.905 1.585 ;
        RECT  6.745 2.505 6.905 2.765 ;
        RECT  6.690 0.455 6.890 0.715 ;
        RECT  6.550 1.015 6.710 1.585 ;
        RECT  6.270 1.795 6.635 2.055 ;
        RECT  6.310 1.015 6.550 1.175 ;
        RECT  6.130 1.380 6.270 2.225 ;
        RECT  6.110 0.995 6.130 2.225 ;
        RECT  5.970 0.995 6.110 1.540 ;
        RECT  6.100 2.065 6.110 2.225 ;
        RECT  5.840 2.065 6.100 2.325 ;
        RECT  5.935 2.520 6.095 3.105 ;
        RECT  5.560 0.995 5.970 1.155 ;
        RECT  3.915 2.520 5.935 2.680 ;
        RECT  5.300 0.895 5.560 1.155 ;
        RECT  4.550 2.860 4.810 3.120 ;
        RECT  4.255 2.170 4.680 2.330 ;
        RECT  3.575 2.860 4.550 3.020 ;
        RECT  4.095 2.015 4.255 2.330 ;
        RECT  3.940 1.045 4.110 1.305 ;
        RECT  3.940 2.015 4.095 2.175 ;
        RECT  3.780 1.045 3.940 2.175 ;
        RECT  3.755 2.355 3.915 2.680 ;
        RECT  3.585 1.575 3.780 1.835 ;
        RECT  2.555 2.355 3.755 2.515 ;
        RECT  3.340 1.045 3.600 1.305 ;
        RECT  3.120 2.015 3.595 2.175 ;
        RECT  3.415 2.695 3.575 3.020 ;
        RECT  2.895 2.695 3.415 2.855 ;
        RECT  3.120 1.095 3.340 1.305 ;
        RECT  2.960 1.095 3.120 2.175 ;
        RECT  2.615 1.095 2.960 1.255 ;
        RECT  2.735 2.695 2.895 3.135 ;
        RECT  1.365 2.975 2.735 3.135 ;
        RECT  2.455 0.835 2.615 1.255 ;
        RECT  2.395 2.355 2.555 2.735 ;
        RECT  2.115 0.835 2.455 0.995 ;
        RECT  1.705 2.575 2.395 2.735 ;
        RECT  2.115 1.175 2.275 1.335 ;
        RECT  2.115 2.130 2.215 2.390 ;
        RECT  1.855 0.770 2.115 0.995 ;
        RECT  1.955 1.175 2.115 2.390 ;
        RECT  1.705 1.210 1.725 1.470 ;
        RECT  1.545 1.210 1.705 2.735 ;
        RECT  1.515 1.210 1.545 2.390 ;
        RECT  1.465 1.210 1.515 1.470 ;
        RECT  1.445 2.130 1.515 2.390 ;
        RECT  1.205 2.580 1.365 3.135 ;
        RECT  0.385 2.580 1.205 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.115 1.025 0.225 2.515 ;
    END
END SMDFFHQX2

MACRO SMDFFHQX1
    CLASS CORE ;
    FOREIGN SMDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.360 1.385 4.900 1.545 ;
        RECT  4.200 0.585 4.360 1.545 ;
        RECT  2.955 0.585 4.200 0.745 ;
        RECT  2.795 0.470 2.955 0.745 ;
        RECT  2.460 0.470 2.795 0.630 ;
        RECT  2.300 0.465 2.460 0.630 ;
        RECT  1.645 0.465 2.300 0.625 ;
        RECT  1.485 0.465 1.645 0.805 ;
        RECT  1.305 0.645 1.485 0.805 ;
        RECT  1.145 0.645 1.305 1.380 ;
        RECT  1.045 1.105 1.145 1.380 ;
        RECT  0.795 1.220 1.045 1.380 ;
        RECT  0.770 1.220 0.795 1.580 ;
        RECT  0.715 1.220 0.770 1.680 ;
        RECT  0.610 1.220 0.715 1.730 ;
        RECT  0.585 1.290 0.610 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.725 5.380 1.885 ;
        RECT  3.975 1.700 4.015 1.990 ;
        RECT  3.815 1.660 3.975 1.990 ;
        RECT  3.805 1.700 3.815 1.990 ;
        END
        ANTENNAGATEAREA     0.0975 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.025 1.105 14.135 2.175 ;
        RECT  13.865 0.695 14.025 2.680 ;
        RECT  13.565 0.695 13.865 0.855 ;
        RECT  13.675 2.520 13.865 2.680 ;
        RECT  13.505 2.520 13.675 2.995 ;
        RECT  13.305 0.595 13.565 0.855 ;
        RECT  13.245 2.520 13.505 3.165 ;
        END
        ANTENNADIFFAREA     0.3808 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.535 2.635 1.990 ;
        RECT  2.305 1.535 2.425 1.895 ;
        END
        ANTENNAGATEAREA     0.0923 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.040 0.880 7.235 1.620 ;
        RECT  7.025 0.880 7.040 1.170 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  7.755 1.290 8.155 1.620 ;
        END
        ANTENNAGATEAREA     0.1261 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.025 -0.250 14.260 0.250 ;
        RECT  12.765 -0.250 13.025 0.405 ;
        RECT  10.970 -0.250 12.765 0.250 ;
        RECT  10.710 -0.250 10.970 0.405 ;
        RECT  9.290 -0.250 10.710 0.250 ;
        RECT  9.030 -0.250 9.290 0.405 ;
        RECT  7.340 -0.250 9.030 0.250 ;
        RECT  7.080 -0.250 7.340 0.405 ;
        RECT  5.530 -0.250 7.080 0.250 ;
        RECT  5.270 -0.250 5.530 0.405 ;
        RECT  4.515 -0.250 5.270 0.250 ;
        RECT  4.255 -0.250 4.515 0.405 ;
        RECT  3.395 -0.250 4.255 0.250 ;
        RECT  3.135 -0.250 3.395 0.405 ;
        RECT  0.815 -0.250 3.135 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.985 3.440 14.260 3.940 ;
        RECT  12.725 2.615 12.985 3.940 ;
        RECT  11.160 3.440 12.725 3.940 ;
        RECT  10.900 3.285 11.160 3.940 ;
        RECT  9.400 3.440 10.900 3.940 ;
        RECT  9.140 3.285 9.400 3.940 ;
        RECT  7.480 3.440 9.140 3.940 ;
        RECT  7.220 3.285 7.480 3.940 ;
        RECT  5.540 3.440 7.220 3.940 ;
        RECT  5.280 3.285 5.540 3.940 ;
        RECT  4.775 3.440 5.280 3.940 ;
        RECT  4.515 2.925 4.775 3.940 ;
        RECT  3.765 3.440 4.515 3.940 ;
        RECT  3.505 3.285 3.765 3.940 ;
        RECT  2.615 3.440 3.505 3.940 ;
        RECT  2.355 3.115 2.615 3.940 ;
        RECT  0.815 3.440 2.355 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.535 1.105 13.645 2.165 ;
        RECT  13.485 1.105 13.535 2.285 ;
        RECT  13.385 1.105 13.485 1.365 ;
        RECT  13.275 2.005 13.485 2.285 ;
        RECT  13.205 1.560 13.305 1.820 ;
        RECT  12.725 2.005 13.275 2.165 ;
        RECT  13.045 1.310 13.205 1.820 ;
        RECT  12.725 1.310 13.045 1.470 ;
        RECT  12.565 0.745 12.725 1.470 ;
        RECT  12.565 1.785 12.725 2.165 ;
        RECT  12.045 0.745 12.565 0.905 ;
        RECT  12.225 1.085 12.385 3.215 ;
        RECT  11.595 3.055 12.225 3.215 ;
        RECT  11.885 0.745 12.045 2.795 ;
        RECT  11.770 0.975 11.885 1.235 ;
        RECT  11.640 0.570 11.690 0.730 ;
        RECT  11.430 0.570 11.640 0.745 ;
        RECT  11.435 2.940 11.595 3.215 ;
        RECT  11.560 2.135 11.585 2.760 ;
        RECT  11.400 1.035 11.560 2.760 ;
        RECT  10.280 2.940 11.435 3.100 ;
        RECT  8.850 0.585 11.430 0.745 ;
        RECT  11.260 1.035 11.400 1.295 ;
        RECT  11.325 2.135 11.400 2.760 ;
        RECT  10.530 2.600 11.325 2.760 ;
        RECT  10.785 1.635 11.220 1.895 ;
        RECT  10.625 1.025 10.785 2.420 ;
        RECT  10.180 1.025 10.625 1.185 ;
        RECT  9.850 2.260 10.625 2.420 ;
        RECT  9.845 1.635 10.310 1.895 ;
        RECT  10.120 2.605 10.280 3.100 ;
        RECT  10.020 0.925 10.180 1.185 ;
        RECT  9.670 2.605 10.120 2.765 ;
        RECT  8.755 2.945 9.940 3.105 ;
        RECT  9.840 1.635 9.845 2.065 ;
        RECT  9.680 1.135 9.840 2.065 ;
        RECT  9.450 1.135 9.680 1.295 ;
        RECT  9.670 1.905 9.680 2.065 ;
        RECT  9.510 1.905 9.670 2.765 ;
        RECT  8.340 2.605 9.510 2.765 ;
        RECT  8.850 1.565 9.500 1.725 ;
        RECT  9.290 1.035 9.450 1.295 ;
        RECT  8.710 0.585 8.850 2.405 ;
        RECT  8.595 2.945 8.755 3.135 ;
        RECT  8.690 0.510 8.710 2.405 ;
        RECT  8.450 0.510 8.690 0.770 ;
        RECT  7.910 2.245 8.690 2.405 ;
        RECT  7.820 2.975 8.595 3.135 ;
        RECT  8.335 0.950 8.495 2.035 ;
        RECT  8.080 2.605 8.340 2.775 ;
        RECT  8.270 0.950 8.335 1.110 ;
        RECT  7.800 1.875 8.335 2.035 ;
        RECT  8.110 0.440 8.270 1.110 ;
        RECT  7.670 0.440 8.110 0.600 ;
        RECT  7.575 2.605 8.080 2.765 ;
        RECT  7.575 0.950 7.930 1.110 ;
        RECT  7.660 2.945 7.820 3.135 ;
        RECT  6.520 2.945 7.660 3.105 ;
        RECT  7.415 0.950 7.575 2.765 ;
        RECT  6.860 2.170 7.080 2.430 ;
        RECT  6.845 1.350 6.860 2.430 ;
        RECT  6.820 0.905 6.845 2.430 ;
        RECT  6.700 0.905 6.820 2.380 ;
        RECT  6.685 0.905 6.700 1.510 ;
        RECT  6.505 2.140 6.520 3.105 ;
        RECT  6.345 0.545 6.505 3.105 ;
        RECT  6.325 0.545 6.345 0.705 ;
        RECT  5.115 2.945 6.345 3.105 ;
        RECT  6.065 0.445 6.325 0.705 ;
        RECT  6.060 1.015 6.150 2.715 ;
        RECT  5.990 1.015 6.060 2.765 ;
        RECT  5.850 1.015 5.990 1.175 ;
        RECT  5.960 1.850 5.990 2.110 ;
        RECT  5.800 2.505 5.990 2.765 ;
        RECT  5.720 1.370 5.810 1.630 ;
        RECT  5.670 1.370 5.720 2.225 ;
        RECT  5.560 1.045 5.670 2.225 ;
        RECT  5.510 1.045 5.560 1.540 ;
        RECT  5.485 2.065 5.560 2.225 ;
        RECT  5.100 1.045 5.510 1.205 ;
        RECT  5.225 2.065 5.485 2.325 ;
        RECT  4.955 2.510 5.115 3.105 ;
        RECT  4.840 0.945 5.100 1.205 ;
        RECT  3.295 2.510 4.955 2.670 ;
        RECT  4.075 2.850 4.335 3.110 ;
        RECT  3.625 2.170 4.195 2.330 ;
        RECT  2.955 2.850 4.075 3.010 ;
        RECT  3.625 0.965 3.765 1.225 ;
        RECT  3.465 0.965 3.625 2.330 ;
        RECT  3.155 1.635 3.465 1.895 ;
        RECT  3.135 2.435 3.295 2.670 ;
        RECT  2.975 1.125 3.255 1.385 ;
        RECT  2.975 2.095 3.255 2.255 ;
        RECT  1.705 2.435 3.135 2.595 ;
        RECT  2.815 1.125 2.975 2.255 ;
        RECT  2.795 2.775 2.955 3.010 ;
        RECT  2.615 1.125 2.815 1.285 ;
        RECT  1.365 2.775 2.795 2.935 ;
        RECT  2.455 0.810 2.615 1.285 ;
        RECT  2.105 0.810 2.455 0.970 ;
        RECT  2.115 1.175 2.275 1.335 ;
        RECT  2.115 2.095 2.215 2.255 ;
        RECT  1.955 1.175 2.115 2.255 ;
        RECT  1.845 0.805 2.105 0.970 ;
        RECT  1.675 2.150 1.705 2.595 ;
        RECT  1.545 1.035 1.675 2.595 ;
        RECT  1.515 1.035 1.545 2.410 ;
        RECT  1.445 2.150 1.515 2.410 ;
        RECT  1.205 2.580 1.365 2.935 ;
        RECT  0.385 2.580 1.205 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.125 1.025 0.225 2.520 ;
        RECT  0.115 1.035 0.125 2.520 ;
    END
END SMDFFHQX1

MACRO SEDFFHQX8
    CLASS CORE ;
    FOREIGN SEDFFHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.620 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.990 1.255 2.400 ;
        RECT  0.975 1.565 1.235 2.400 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.335 6.305 1.495 ;
        RECT  5.740 1.105 5.855 1.495 ;
        RECT  5.580 0.650 5.740 1.495 ;
        RECT  4.415 0.650 5.580 0.810 ;
        RECT  4.255 0.470 4.415 0.810 ;
        RECT  1.505 0.470 4.255 0.630 ;
        RECT  1.435 0.430 1.505 0.630 ;
        RECT  1.230 0.430 1.435 0.745 ;
        RECT  0.795 0.585 1.230 0.745 ;
        RECT  0.715 0.585 0.795 1.680 ;
        RECT  0.635 0.585 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.955 1.515 21.035 1.765 ;
        RECT  20.695 0.695 20.955 2.895 ;
        RECT  19.930 1.290 20.695 1.990 ;
        RECT  19.670 0.695 19.930 2.920 ;
        END
        ANTENNADIFFAREA     1.5960 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.725 6.770 1.885 ;
        RECT  5.645 1.700 5.855 1.990 ;
        RECT  5.335 1.700 5.645 1.860 ;
        RECT  5.175 1.575 5.335 1.860 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.670 2.805 2.030 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.975 1.290 9.995 1.580 ;
        RECT  9.815 1.155 9.975 1.580 ;
        RECT  9.585 1.290 9.815 1.580 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.465 -0.250 21.620 0.250 ;
        RECT  21.205 -0.250 21.465 1.115 ;
        RECT  20.440 -0.250 21.205 0.250 ;
        RECT  20.180 -0.250 20.440 0.940 ;
        RECT  19.415 -0.250 20.180 0.250 ;
        RECT  19.155 -0.250 19.415 1.295 ;
        RECT  18.630 -0.250 19.155 0.250 ;
        RECT  18.370 -0.250 18.630 0.405 ;
        RECT  9.835 -0.250 18.370 0.250 ;
        RECT  9.575 -0.250 9.835 0.405 ;
        RECT  8.785 -0.250 9.575 0.250 ;
        RECT  8.525 -0.250 8.785 0.405 ;
        RECT  7.095 -0.250 8.525 0.250 ;
        RECT  6.835 -0.250 7.095 0.405 ;
        RECT  6.075 -0.250 6.835 0.250 ;
        RECT  5.815 -0.250 6.075 0.405 ;
        RECT  4.855 -0.250 5.815 0.250 ;
        RECT  4.595 -0.250 4.855 0.405 ;
        RECT  0.815 -0.250 4.595 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.465 3.440 21.620 3.940 ;
        RECT  21.205 2.255 21.465 3.940 ;
        RECT  20.440 3.440 21.205 3.940 ;
        RECT  20.180 2.255 20.440 3.940 ;
        RECT  19.385 3.440 20.180 3.940 ;
        RECT  19.125 3.285 19.385 3.940 ;
        RECT  18.505 3.440 19.125 3.940 ;
        RECT  18.245 3.285 18.505 3.940 ;
        RECT  15.910 3.440 18.245 3.940 ;
        RECT  15.650 3.285 15.910 3.940 ;
        RECT  14.795 3.440 15.650 3.940 ;
        RECT  14.535 3.285 14.795 3.940 ;
        RECT  13.520 3.440 14.535 3.940 ;
        RECT  13.260 3.285 13.520 3.940 ;
        RECT  11.790 3.440 13.260 3.940 ;
        RECT  11.530 3.285 11.790 3.940 ;
        RECT  10.710 3.440 11.530 3.940 ;
        RECT  10.450 3.285 10.710 3.940 ;
        RECT  8.725 3.440 10.450 3.940 ;
        RECT  8.465 3.285 8.725 3.940 ;
        RECT  6.965 3.440 8.465 3.940 ;
        RECT  6.705 3.285 6.965 3.940 ;
        RECT  6.110 3.440 6.705 3.940 ;
        RECT  5.850 2.945 6.110 3.940 ;
        RECT  5.100 3.440 5.850 3.940 ;
        RECT  4.840 3.285 5.100 3.940 ;
        RECT  4.360 3.405 4.840 3.940 ;
        RECT  4.100 3.095 4.360 3.940 ;
        RECT  0.870 3.440 4.100 3.940 ;
        RECT  0.610 2.925 0.870 3.940 ;
        RECT  0.000 3.440 0.610 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.895 2.575 18.935 2.835 ;
        RECT  18.735 0.845 18.895 2.835 ;
        RECT  18.625 0.845 18.735 1.225 ;
        RECT  18.640 1.885 18.735 2.145 ;
        RECT  18.675 2.575 18.735 2.835 ;
        RECT  18.190 0.845 18.625 1.005 ;
        RECT  18.445 1.405 18.555 1.665 ;
        RECT  18.285 1.185 18.445 2.880 ;
        RECT  17.850 1.185 18.285 1.345 ;
        RECT  16.820 2.720 18.285 2.880 ;
        RECT  18.030 0.470 18.190 1.005 ;
        RECT  17.945 1.530 18.105 2.535 ;
        RECT  14.490 0.470 18.030 0.630 ;
        RECT  17.510 1.530 17.945 1.690 ;
        RECT  17.360 2.375 17.945 2.535 ;
        RECT  17.690 0.910 17.850 1.345 ;
        RECT  17.605 1.875 17.765 2.190 ;
        RECT  17.360 0.910 17.690 1.070 ;
        RECT  17.170 1.875 17.605 2.035 ;
        RECT  17.335 3.060 17.595 3.260 ;
        RECT  17.350 1.250 17.510 1.690 ;
        RECT  17.100 0.810 17.360 1.070 ;
        RECT  17.200 2.220 17.360 2.535 ;
        RECT  16.820 1.250 17.350 1.410 ;
        RECT  16.250 3.060 17.335 3.220 ;
        RECT  16.820 2.220 17.200 2.380 ;
        RECT  17.010 1.635 17.170 2.035 ;
        RECT  16.230 0.810 17.100 0.970 ;
        RECT  15.540 1.635 17.010 1.795 ;
        RECT  16.560 1.155 16.820 1.410 ;
        RECT  16.560 2.120 16.820 2.380 ;
        RECT  16.660 2.565 16.820 2.880 ;
        RECT  16.280 2.565 16.660 2.725 ;
        RECT  15.880 1.250 16.560 1.410 ;
        RECT  15.370 2.120 16.560 2.280 ;
        RECT  16.020 2.465 16.280 2.725 ;
        RECT  16.090 2.940 16.250 3.220 ;
        RECT  16.070 0.810 16.230 1.070 ;
        RECT  14.160 2.940 16.090 3.100 ;
        RECT  15.720 0.910 15.880 1.410 ;
        RECT  15.370 0.910 15.720 1.070 ;
        RECT  15.380 1.250 15.540 1.795 ;
        RECT  14.760 1.250 15.380 1.410 ;
        RECT  15.110 0.810 15.370 1.070 ;
        RECT  15.110 2.120 15.370 2.760 ;
        RECT  14.940 1.635 15.200 1.850 ;
        RECT  14.340 2.600 15.110 2.760 ;
        RECT  13.955 1.690 14.940 1.850 ;
        RECT  14.600 0.810 14.760 1.410 ;
        RECT  14.145 0.810 14.600 0.970 ;
        RECT  14.330 0.430 14.490 0.630 ;
        RECT  13.695 0.430 14.330 0.590 ;
        RECT  14.000 2.605 14.160 3.100 ;
        RECT  13.885 0.770 14.145 0.970 ;
        RECT  12.195 2.605 14.000 2.765 ;
        RECT  13.875 1.150 13.955 2.320 ;
        RECT  11.425 0.810 13.885 0.970 ;
        RECT  13.795 1.150 13.875 2.425 ;
        RECT  12.435 1.150 13.795 1.310 ;
        RECT  13.615 2.160 13.795 2.425 ;
        RECT  13.535 0.430 13.695 0.630 ;
        RECT  12.200 1.680 13.615 1.840 ;
        RECT  12.655 2.160 13.615 2.320 ;
        RECT  10.355 0.470 13.535 0.630 ;
        RECT  12.225 2.945 12.825 3.215 ;
        RECT  12.395 2.160 12.655 2.420 ;
        RECT  7.930 2.945 12.225 3.105 ;
        RECT  12.195 1.195 12.200 1.840 ;
        RECT  12.035 1.195 12.195 2.765 ;
        RECT  11.755 1.195 12.035 1.355 ;
        RECT  8.270 2.605 12.035 2.765 ;
        RECT  11.425 1.610 11.850 1.885 ;
        RECT  11.265 0.810 11.425 2.325 ;
        RECT  10.760 1.125 11.265 1.385 ;
        RECT  11.250 2.165 11.265 2.325 ;
        RECT  10.990 2.165 11.250 2.425 ;
        RECT  10.370 1.650 11.080 1.910 ;
        RECT  9.905 2.265 10.990 2.425 ;
        RECT  10.370 0.925 10.415 1.085 ;
        RECT  10.210 0.925 10.370 1.995 ;
        RECT  10.195 0.470 10.355 0.745 ;
        RECT  10.155 0.925 10.210 1.085 ;
        RECT  9.430 1.835 10.210 1.995 ;
        RECT  9.585 0.585 10.195 0.745 ;
        RECT  9.645 2.210 9.905 2.425 ;
        RECT  9.425 0.585 9.585 1.100 ;
        RECT  9.170 1.735 9.430 1.995 ;
        RECT  8.710 0.940 9.425 1.100 ;
        RECT  9.085 0.500 9.245 0.760 ;
        RECT  8.270 0.600 9.085 0.760 ;
        RECT  8.450 0.940 8.710 1.245 ;
        RECT  8.110 0.600 8.270 2.765 ;
        RECT  7.770 0.495 7.930 3.105 ;
        RECT  7.625 0.495 7.770 0.755 ;
        RECT  6.450 2.945 7.770 3.105 ;
        RECT  7.575 1.005 7.590 2.155 ;
        RECT  7.455 1.005 7.575 2.190 ;
        RECT  7.430 1.005 7.455 2.740 ;
        RECT  7.315 1.005 7.430 1.265 ;
        RECT  7.295 1.895 7.430 2.740 ;
        RECT  7.145 2.580 7.295 2.740 ;
        RECT  7.110 1.450 7.250 1.710 ;
        RECT  6.950 0.995 7.110 2.225 ;
        RECT  6.510 0.995 6.950 1.155 ;
        RECT  6.775 2.065 6.950 2.225 ;
        RECT  6.615 2.065 6.775 2.325 ;
        RECT  6.250 0.895 6.510 1.155 ;
        RECT  6.290 2.510 6.450 3.105 ;
        RECT  5.080 2.510 6.290 2.670 ;
        RECT  4.700 2.860 5.670 3.020 ;
        RECT  5.460 2.170 5.530 2.330 ;
        RECT  5.270 2.075 5.460 2.330 ;
        RECT  4.965 2.075 5.270 2.235 ;
        RECT  4.965 1.045 5.185 1.305 ;
        RECT  4.920 2.415 5.080 2.670 ;
        RECT  4.925 1.045 4.965 2.235 ;
        RECT  4.805 1.145 4.925 2.235 ;
        RECT  3.580 2.415 4.920 2.575 ;
        RECT  4.460 1.635 4.805 1.895 ;
        RECT  4.540 2.755 4.700 3.020 ;
        RECT  4.075 1.025 4.625 1.285 ;
        RECT  3.920 2.755 4.540 2.915 ;
        RECT  4.075 2.075 4.520 2.235 ;
        RECT  3.915 0.810 4.075 2.235 ;
        RECT  3.760 2.755 3.920 3.220 ;
        RECT  1.815 0.810 3.915 0.970 ;
        RECT  1.250 3.060 3.760 3.220 ;
        RECT  3.580 1.155 3.735 1.315 ;
        RECT  3.420 1.155 3.580 2.820 ;
        RECT  1.730 2.660 3.420 2.820 ;
        RECT  2.985 1.250 3.145 2.480 ;
        RECT  2.240 2.220 2.985 2.380 ;
        RECT  2.240 1.250 2.245 1.510 ;
        RECT  2.080 1.250 2.240 2.480 ;
        RECT  1.985 1.250 2.080 1.510 ;
        RECT  1.980 2.220 2.080 2.480 ;
        RECT  1.730 1.170 1.735 1.430 ;
        RECT  1.570 1.170 1.730 2.820 ;
        RECT  1.475 1.170 1.570 1.430 ;
        RECT  1.470 2.420 1.570 2.680 ;
        RECT  1.090 2.580 1.250 3.220 ;
        RECT  0.385 2.580 1.090 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.115 1.025 0.225 2.520 ;
    END
END SEDFFHQX8

MACRO SEDFFHQX4
    CLASS CORE ;
    FOREIGN SEDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.700 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.990 1.255 2.400 ;
        RECT  0.975 1.565 1.235 2.400 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.335 6.305 1.495 ;
        RECT  5.740 1.105 5.855 1.495 ;
        RECT  5.580 0.650 5.740 1.495 ;
        RECT  4.415 0.650 5.580 0.810 ;
        RECT  4.255 0.470 4.415 0.810 ;
        RECT  1.505 0.470 4.255 0.630 ;
        RECT  1.435 0.430 1.505 0.630 ;
        RECT  1.230 0.430 1.435 0.745 ;
        RECT  0.795 0.585 1.230 0.745 ;
        RECT  0.715 0.585 0.795 1.680 ;
        RECT  0.635 0.585 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.930 1.515 20.115 1.765 ;
        RECT  19.670 0.695 19.930 2.920 ;
        RECT  19.595 1.695 19.670 2.400 ;
        RECT  19.445 1.700 19.595 2.400 ;
        END
        ANTENNADIFFAREA     0.7980 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.725 6.770 1.885 ;
        RECT  5.645 1.700 5.855 1.990 ;
        RECT  5.335 1.700 5.645 1.860 ;
        RECT  5.175 1.575 5.335 1.860 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.670 2.805 2.030 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.975 1.290 9.995 1.580 ;
        RECT  9.815 1.155 9.975 1.580 ;
        RECT  9.585 1.290 9.815 1.580 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.440 -0.250 20.700 0.250 ;
        RECT  20.180 -0.250 20.440 1.115 ;
        RECT  19.415 -0.250 20.180 0.250 ;
        RECT  19.155 -0.250 19.415 1.295 ;
        RECT  18.630 -0.250 19.155 0.250 ;
        RECT  18.370 -0.250 18.630 0.405 ;
        RECT  9.835 -0.250 18.370 0.250 ;
        RECT  9.575 -0.250 9.835 0.405 ;
        RECT  8.785 -0.250 9.575 0.250 ;
        RECT  8.525 -0.250 8.785 0.405 ;
        RECT  7.095 -0.250 8.525 0.250 ;
        RECT  6.835 -0.250 7.095 0.405 ;
        RECT  6.075 -0.250 6.835 0.250 ;
        RECT  5.815 -0.250 6.075 0.405 ;
        RECT  4.855 -0.250 5.815 0.250 ;
        RECT  4.595 -0.250 4.855 0.405 ;
        RECT  0.815 -0.250 4.595 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.440 3.440 20.700 3.940 ;
        RECT  20.180 2.255 20.440 3.940 ;
        RECT  19.385 3.440 20.180 3.940 ;
        RECT  19.125 3.285 19.385 3.940 ;
        RECT  18.505 3.440 19.125 3.940 ;
        RECT  18.245 3.285 18.505 3.940 ;
        RECT  15.910 3.440 18.245 3.940 ;
        RECT  15.650 3.285 15.910 3.940 ;
        RECT  14.795 3.440 15.650 3.940 ;
        RECT  14.535 3.285 14.795 3.940 ;
        RECT  13.520 3.440 14.535 3.940 ;
        RECT  13.260 3.285 13.520 3.940 ;
        RECT  11.790 3.440 13.260 3.940 ;
        RECT  11.530 3.285 11.790 3.940 ;
        RECT  10.710 3.440 11.530 3.940 ;
        RECT  10.450 3.285 10.710 3.940 ;
        RECT  8.725 3.440 10.450 3.940 ;
        RECT  8.465 3.285 8.725 3.940 ;
        RECT  6.965 3.440 8.465 3.940 ;
        RECT  6.705 3.285 6.965 3.940 ;
        RECT  6.110 3.440 6.705 3.940 ;
        RECT  5.850 2.945 6.110 3.940 ;
        RECT  5.100 3.440 5.850 3.940 ;
        RECT  4.840 3.285 5.100 3.940 ;
        RECT  4.360 3.405 4.840 3.940 ;
        RECT  4.100 3.095 4.360 3.940 ;
        RECT  0.870 3.440 4.100 3.940 ;
        RECT  0.610 2.925 0.870 3.940 ;
        RECT  0.000 3.440 0.610 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.895 2.575 18.935 2.835 ;
        RECT  18.735 0.845 18.895 2.835 ;
        RECT  18.625 0.845 18.735 1.225 ;
        RECT  18.640 1.885 18.735 2.145 ;
        RECT  18.675 2.575 18.735 2.835 ;
        RECT  18.190 0.845 18.625 1.005 ;
        RECT  18.445 1.405 18.555 1.665 ;
        RECT  18.285 1.185 18.445 2.880 ;
        RECT  17.850 1.185 18.285 1.345 ;
        RECT  16.820 2.720 18.285 2.880 ;
        RECT  18.030 0.470 18.190 1.005 ;
        RECT  17.945 1.530 18.105 2.535 ;
        RECT  14.490 0.470 18.030 0.630 ;
        RECT  17.510 1.530 17.945 1.690 ;
        RECT  17.360 2.375 17.945 2.535 ;
        RECT  17.690 0.910 17.850 1.345 ;
        RECT  17.605 1.875 17.765 2.190 ;
        RECT  17.360 0.910 17.690 1.070 ;
        RECT  17.170 1.875 17.605 2.035 ;
        RECT  17.335 3.060 17.595 3.260 ;
        RECT  17.350 1.250 17.510 1.690 ;
        RECT  17.100 0.810 17.360 1.070 ;
        RECT  17.200 2.220 17.360 2.535 ;
        RECT  16.820 1.250 17.350 1.410 ;
        RECT  16.250 3.060 17.335 3.220 ;
        RECT  16.820 2.220 17.200 2.380 ;
        RECT  17.010 1.635 17.170 2.035 ;
        RECT  16.230 0.810 17.100 0.970 ;
        RECT  15.540 1.635 17.010 1.795 ;
        RECT  16.560 1.155 16.820 1.410 ;
        RECT  16.560 2.120 16.820 2.380 ;
        RECT  16.660 2.565 16.820 2.880 ;
        RECT  16.280 2.565 16.660 2.725 ;
        RECT  15.880 1.250 16.560 1.410 ;
        RECT  15.370 2.120 16.560 2.280 ;
        RECT  16.020 2.465 16.280 2.725 ;
        RECT  16.090 2.940 16.250 3.220 ;
        RECT  16.070 0.810 16.230 1.070 ;
        RECT  14.160 2.940 16.090 3.100 ;
        RECT  15.720 0.910 15.880 1.410 ;
        RECT  15.370 0.910 15.720 1.070 ;
        RECT  15.380 1.250 15.540 1.795 ;
        RECT  14.760 1.250 15.380 1.410 ;
        RECT  15.110 0.810 15.370 1.070 ;
        RECT  15.110 2.120 15.370 2.760 ;
        RECT  14.940 1.635 15.200 1.850 ;
        RECT  14.340 2.600 15.110 2.760 ;
        RECT  13.955 1.690 14.940 1.850 ;
        RECT  14.600 0.810 14.760 1.410 ;
        RECT  14.145 0.810 14.600 0.970 ;
        RECT  14.330 0.430 14.490 0.630 ;
        RECT  13.695 0.430 14.330 0.590 ;
        RECT  14.000 2.605 14.160 3.100 ;
        RECT  13.885 0.770 14.145 0.970 ;
        RECT  12.195 2.605 14.000 2.765 ;
        RECT  13.875 1.150 13.955 2.320 ;
        RECT  11.425 0.810 13.885 0.970 ;
        RECT  13.795 1.150 13.875 2.425 ;
        RECT  12.435 1.150 13.795 1.310 ;
        RECT  13.615 2.160 13.795 2.425 ;
        RECT  13.535 0.430 13.695 0.630 ;
        RECT  12.200 1.680 13.615 1.840 ;
        RECT  12.655 2.160 13.615 2.320 ;
        RECT  10.355 0.470 13.535 0.630 ;
        RECT  12.225 2.945 12.825 3.215 ;
        RECT  12.395 2.160 12.655 2.420 ;
        RECT  7.930 2.945 12.225 3.105 ;
        RECT  12.195 1.195 12.200 1.840 ;
        RECT  12.035 1.195 12.195 2.765 ;
        RECT  11.755 1.195 12.035 1.355 ;
        RECT  8.270 2.605 12.035 2.765 ;
        RECT  11.425 1.610 11.850 1.885 ;
        RECT  11.265 0.810 11.425 2.325 ;
        RECT  10.760 1.125 11.265 1.385 ;
        RECT  11.250 2.165 11.265 2.325 ;
        RECT  10.990 2.165 11.250 2.425 ;
        RECT  10.370 1.650 11.080 1.910 ;
        RECT  9.905 2.265 10.990 2.425 ;
        RECT  10.370 0.925 10.415 1.085 ;
        RECT  10.210 0.925 10.370 1.995 ;
        RECT  10.195 0.470 10.355 0.745 ;
        RECT  10.155 0.925 10.210 1.085 ;
        RECT  9.430 1.835 10.210 1.995 ;
        RECT  9.585 0.585 10.195 0.745 ;
        RECT  9.645 2.210 9.905 2.425 ;
        RECT  9.425 0.585 9.585 1.100 ;
        RECT  9.170 1.735 9.430 1.995 ;
        RECT  8.710 0.940 9.425 1.100 ;
        RECT  9.085 0.500 9.245 0.760 ;
        RECT  8.270 0.600 9.085 0.760 ;
        RECT  8.450 0.940 8.710 1.245 ;
        RECT  8.110 0.600 8.270 2.765 ;
        RECT  7.770 0.495 7.930 3.105 ;
        RECT  7.625 0.495 7.770 0.755 ;
        RECT  6.450 2.945 7.770 3.105 ;
        RECT  7.575 1.005 7.590 2.155 ;
        RECT  7.455 1.005 7.575 2.190 ;
        RECT  7.430 1.005 7.455 2.740 ;
        RECT  7.315 1.005 7.430 1.265 ;
        RECT  7.295 1.895 7.430 2.740 ;
        RECT  7.145 2.580 7.295 2.740 ;
        RECT  7.110 1.450 7.250 1.710 ;
        RECT  6.950 0.995 7.110 2.225 ;
        RECT  6.510 0.995 6.950 1.155 ;
        RECT  6.775 2.065 6.950 2.225 ;
        RECT  6.615 2.065 6.775 2.325 ;
        RECT  6.250 0.895 6.510 1.155 ;
        RECT  6.290 2.510 6.450 3.105 ;
        RECT  5.080 2.510 6.290 2.670 ;
        RECT  4.700 2.860 5.670 3.020 ;
        RECT  5.460 2.170 5.530 2.330 ;
        RECT  5.270 2.075 5.460 2.330 ;
        RECT  4.965 2.075 5.270 2.235 ;
        RECT  4.965 1.045 5.185 1.305 ;
        RECT  4.920 2.415 5.080 2.670 ;
        RECT  4.925 1.045 4.965 2.235 ;
        RECT  4.805 1.145 4.925 2.235 ;
        RECT  3.580 2.415 4.920 2.575 ;
        RECT  4.460 1.635 4.805 1.895 ;
        RECT  4.540 2.755 4.700 3.020 ;
        RECT  4.075 1.025 4.625 1.285 ;
        RECT  3.920 2.755 4.540 2.915 ;
        RECT  4.075 2.075 4.520 2.235 ;
        RECT  3.915 0.810 4.075 2.235 ;
        RECT  3.760 2.755 3.920 3.220 ;
        RECT  1.815 0.810 3.915 0.970 ;
        RECT  1.250 3.060 3.760 3.220 ;
        RECT  3.580 1.155 3.735 1.315 ;
        RECT  3.420 1.155 3.580 2.820 ;
        RECT  1.730 2.660 3.420 2.820 ;
        RECT  2.985 1.250 3.145 2.480 ;
        RECT  2.240 2.220 2.985 2.380 ;
        RECT  2.240 1.250 2.245 1.510 ;
        RECT  2.080 1.250 2.240 2.480 ;
        RECT  1.985 1.250 2.080 1.510 ;
        RECT  1.980 2.220 2.080 2.480 ;
        RECT  1.730 1.170 1.735 1.430 ;
        RECT  1.570 1.170 1.730 2.820 ;
        RECT  1.475 1.170 1.570 1.430 ;
        RECT  1.470 2.420 1.570 2.680 ;
        RECT  1.090 2.580 1.250 3.220 ;
        RECT  0.385 2.580 1.090 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.115 1.025 0.225 2.520 ;
    END
END SEDFFHQX4

MACRO SEDFFHQX2
    CLASS CORE ;
    FOREIGN SEDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.100 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.890 1.335 5.255 1.495 ;
        RECT  4.730 1.000 4.890 1.495 ;
        RECT  4.450 1.000 4.730 1.160 ;
        RECT  4.290 0.620 4.450 1.160 ;
        RECT  2.955 0.620 4.290 0.780 ;
        RECT  2.795 0.490 2.955 0.780 ;
        RECT  2.455 0.490 2.795 0.650 ;
        RECT  2.295 0.430 2.455 0.650 ;
        RECT  1.670 0.430 2.295 0.590 ;
        RECT  1.510 0.430 1.670 0.735 ;
        RECT  1.505 0.575 1.510 0.735 ;
        RECT  1.230 0.575 1.505 0.835 ;
        RECT  0.795 0.675 1.230 0.835 ;
        RECT  0.715 0.675 0.795 1.680 ;
        RECT  0.635 0.675 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.860 1.105 15.975 2.585 ;
        RECT  15.820 1.105 15.860 2.895 ;
        RECT  15.660 0.695 15.820 2.895 ;
        RECT  15.560 0.695 15.660 1.295 ;
        RECT  15.600 1.955 15.660 2.895 ;
        RECT  15.305 2.520 15.600 2.810 ;
        END
        ANTENNADIFFAREA     0.7140 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 1.625 5.880 1.885 ;
        RECT  4.935 1.680 5.720 1.840 ;
        RECT  4.930 1.680 4.935 1.990 ;
        RECT  4.725 1.675 4.930 1.990 ;
        RECT  4.285 1.675 4.725 1.835 ;
        RECT  4.125 1.575 4.285 1.835 ;
        END
        ANTENNAGATEAREA     0.1001 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.535 2.635 1.990 ;
        RECT  2.305 1.535 2.425 1.895 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.405 1.285 8.970 1.670 ;
        END
        ANTENNAGATEAREA     0.2327 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.270 -0.250 16.100 0.250 ;
        RECT  14.330 -0.250 15.270 0.405 ;
        RECT  9.010 -0.250 14.330 0.250 ;
        RECT  8.750 -0.250 9.010 0.405 ;
        RECT  7.710 -0.250 8.750 0.250 ;
        RECT  7.450 -0.250 7.710 0.405 ;
        RECT  6.370 -0.250 7.450 0.250 ;
        RECT  5.770 -0.250 6.370 0.405 ;
        RECT  4.880 -0.250 5.770 0.250 ;
        RECT  4.830 -0.250 4.880 0.405 ;
        RECT  4.670 -0.250 4.830 0.795 ;
        RECT  4.620 -0.250 4.670 0.405 ;
        RECT  3.395 -0.250 4.620 0.250 ;
        RECT  3.135 -0.250 3.395 0.405 ;
        RECT  0.815 -0.250 3.135 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.315 3.440 16.100 3.940 ;
        RECT  15.055 3.285 15.315 3.940 ;
        RECT  14.370 3.440 15.055 3.940 ;
        RECT  14.110 2.840 14.370 3.940 ;
        RECT  12.150 3.440 14.110 3.940 ;
        RECT  11.890 3.285 12.150 3.940 ;
        RECT  10.435 3.440 11.890 3.940 ;
        RECT  10.175 3.285 10.435 3.940 ;
        RECT  8.415 3.440 10.175 3.940 ;
        RECT  8.155 3.285 8.415 3.940 ;
        RECT  6.485 3.440 8.155 3.940 ;
        RECT  6.225 3.285 6.485 3.940 ;
        RECT  5.250 3.440 6.225 3.940 ;
        RECT  4.990 2.925 5.250 3.940 ;
        RECT  4.165 3.440 4.990 3.940 ;
        RECT  3.905 3.285 4.165 3.940 ;
        RECT  3.235 3.440 3.905 3.940 ;
        RECT  3.075 3.035 3.235 3.940 ;
        RECT  0.815 3.440 3.075 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.865 2.405 14.950 2.665 ;
        RECT  14.865 0.890 14.890 1.150 ;
        RECT  14.705 0.890 14.865 2.665 ;
        RECT  14.630 0.890 14.705 1.375 ;
        RECT  14.690 2.035 14.705 2.665 ;
        RECT  14.265 2.035 14.690 2.195 ;
        RECT  14.090 1.215 14.630 1.375 ;
        RECT  14.365 1.555 14.525 1.815 ;
        RECT  13.750 1.605 14.365 1.765 ;
        RECT  14.005 2.035 14.265 2.295 ;
        RECT  13.930 0.470 14.090 1.375 ;
        RECT  9.525 0.470 13.930 0.630 ;
        RECT  13.590 0.860 13.750 1.800 ;
        RECT  13.575 2.035 13.735 2.630 ;
        RECT  13.565 3.100 13.615 3.260 ;
        RECT  13.180 0.860 13.590 1.020 ;
        RECT  13.365 1.640 13.590 1.800 ;
        RECT  13.025 2.470 13.575 2.630 ;
        RECT  13.355 2.945 13.565 3.260 ;
        RECT  13.025 1.200 13.410 1.460 ;
        RECT  13.205 1.640 13.365 2.285 ;
        RECT  11.510 2.945 13.355 3.105 ;
        RECT  13.000 1.200 13.025 2.630 ;
        RECT  12.865 0.810 13.000 2.630 ;
        RECT  12.840 0.810 12.865 1.360 ;
        RECT  10.180 0.810 12.840 0.970 ;
        RECT  12.630 2.025 12.685 2.630 ;
        RECT  12.630 1.150 12.660 1.310 ;
        RECT  12.470 1.150 12.630 2.630 ;
        RECT  12.400 1.150 12.470 1.310 ;
        RECT  11.705 2.470 12.470 2.630 ;
        RECT  12.120 1.585 12.290 1.845 ;
        RECT  11.960 1.180 12.120 2.290 ;
        RECT  11.055 1.180 11.960 1.340 ;
        RECT  11.025 2.130 11.960 2.290 ;
        RECT  11.350 2.605 11.510 3.105 ;
        RECT  10.845 1.720 11.485 1.880 ;
        RECT  10.845 2.605 11.350 2.765 ;
        RECT  11.035 3.100 11.115 3.260 ;
        RECT  10.855 2.945 11.035 3.260 ;
        RECT  7.435 2.945 10.855 3.105 ;
        RECT  10.685 1.225 10.845 2.765 ;
        RECT  10.360 1.225 10.685 1.385 ;
        RECT  8.475 2.605 10.685 2.765 ;
        RECT  10.180 1.660 10.505 1.920 ;
        RECT  10.020 0.810 10.180 2.385 ;
        RECT  9.710 0.810 10.020 0.970 ;
        RECT  9.250 2.225 10.020 2.385 ;
        RECT  9.500 1.650 9.825 1.910 ;
        RECT  9.365 0.470 9.525 0.765 ;
        RECT  9.340 0.945 9.500 2.020 ;
        RECT  7.880 0.605 9.365 0.765 ;
        RECT  9.200 0.945 9.340 1.105 ;
        RECT  8.905 1.860 9.340 2.020 ;
        RECT  8.745 1.860 8.905 2.120 ;
        RECT  8.315 1.985 8.475 2.765 ;
        RECT  8.220 0.945 8.345 1.105 ;
        RECT  8.220 1.985 8.315 2.145 ;
        RECT  8.060 0.945 8.220 2.145 ;
        RECT  7.880 2.325 8.135 2.585 ;
        RECT  7.875 0.605 7.880 2.585 ;
        RECT  7.720 0.605 7.875 2.485 ;
        RECT  7.275 1.065 7.435 3.105 ;
        RECT  6.920 1.065 7.275 1.225 ;
        RECT  6.095 2.945 7.275 3.105 ;
        RECT  6.905 1.425 7.065 2.765 ;
        RECT  6.760 0.755 6.920 1.225 ;
        RECT  6.580 1.425 6.905 1.585 ;
        RECT  6.745 2.505 6.905 2.765 ;
        RECT  6.240 1.795 6.635 2.055 ;
        RECT  6.420 0.945 6.580 1.585 ;
        RECT  6.200 0.945 6.420 1.105 ;
        RECT  6.100 1.285 6.240 2.225 ;
        RECT  6.080 1.285 6.100 2.325 ;
        RECT  5.935 2.520 6.095 3.105 ;
        RECT  5.595 1.285 6.080 1.445 ;
        RECT  5.840 2.065 6.080 2.325 ;
        RECT  3.915 2.520 5.935 2.680 ;
        RECT  5.450 0.995 5.595 1.445 ;
        RECT  5.435 0.895 5.450 1.445 ;
        RECT  5.190 0.895 5.435 1.155 ;
        RECT  4.550 2.860 4.810 3.120 ;
        RECT  4.530 2.170 4.680 2.330 ;
        RECT  3.575 2.860 4.550 3.020 ;
        RECT  4.370 2.015 4.530 2.330 ;
        RECT  3.940 2.015 4.370 2.175 ;
        RECT  3.940 1.045 4.110 1.305 ;
        RECT  3.780 1.045 3.940 2.175 ;
        RECT  3.755 2.355 3.915 2.680 ;
        RECT  3.535 1.575 3.780 1.835 ;
        RECT  2.555 2.355 3.755 2.515 ;
        RECT  3.340 1.045 3.600 1.305 ;
        RECT  3.120 2.015 3.595 2.175 ;
        RECT  3.415 2.695 3.575 3.020 ;
        RECT  2.895 2.695 3.415 2.855 ;
        RECT  3.120 1.095 3.340 1.305 ;
        RECT  2.960 1.095 3.120 2.175 ;
        RECT  2.615 1.095 2.960 1.255 ;
        RECT  2.735 2.695 2.895 3.135 ;
        RECT  1.365 2.975 2.735 3.135 ;
        RECT  2.455 0.835 2.615 1.255 ;
        RECT  2.395 2.355 2.555 2.735 ;
        RECT  2.115 0.835 2.455 0.995 ;
        RECT  1.705 2.575 2.395 2.735 ;
        RECT  2.115 1.175 2.275 1.335 ;
        RECT  2.115 2.130 2.215 2.390 ;
        RECT  1.850 0.770 2.115 0.995 ;
        RECT  1.955 1.175 2.115 2.390 ;
        RECT  1.705 1.210 1.725 1.470 ;
        RECT  1.545 1.210 1.705 2.735 ;
        RECT  1.515 1.210 1.545 2.390 ;
        RECT  1.465 1.210 1.515 1.470 ;
        RECT  1.445 2.130 1.515 2.390 ;
        RECT  1.205 2.580 1.365 3.135 ;
        RECT  0.385 2.580 1.205 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.185 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.115 1.025 0.225 2.450 ;
    END
END SEDFFHQX2

MACRO SEDFFHQX1
    CLASS CORE ;
    FOREIGN SEDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.215 1.925 1.255 2.400 ;
        RECT  1.055 1.565 1.215 2.400 ;
        RECT  1.045 1.925 1.055 2.400 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 1.455 4.885 1.615 ;
        RECT  4.420 0.745 4.580 1.615 ;
        RECT  4.265 0.745 4.420 1.355 ;
        RECT  2.975 0.745 4.265 0.905 ;
        RECT  2.815 0.470 2.975 0.905 ;
        RECT  1.530 0.470 2.815 0.630 ;
        RECT  1.230 0.470 1.530 0.805 ;
        RECT  0.795 0.645 1.230 0.805 ;
        RECT  0.665 0.645 0.795 1.580 ;
        RECT  0.610 0.645 0.665 1.730 ;
        RECT  0.585 1.105 0.610 1.730 ;
        RECT  0.505 1.355 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1274 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.540 1.515 14.595 2.585 ;
        RECT  14.395 1.060 14.540 2.810 ;
        RECT  14.380 1.010 14.395 2.810 ;
        RECT  14.235 1.010 14.380 1.270 ;
        RECT  14.220 2.525 14.380 2.810 ;
        RECT  14.135 2.525 14.220 3.170 ;
        RECT  13.960 2.520 14.135 3.170 ;
        RECT  13.925 2.520 13.960 2.995 ;
        END
        ANTENNADIFFAREA     0.5262 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.155 1.675 5.315 1.955 ;
        RECT  4.015 1.795 5.155 1.955 ;
        RECT  3.805 1.700 4.015 2.010 ;
        END
        ANTENNAGATEAREA     0.0975 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.520 2.635 1.990 ;
        RECT  2.295 1.520 2.425 1.920 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.290 7.695 1.905 ;
        END
        ANTENNAGATEAREA     0.1430 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.580 -0.250 14.720 0.250 ;
        RECT  13.320 -0.250 13.580 0.405 ;
        RECT  9.465 -0.250 13.320 0.250 ;
        RECT  9.205 -0.250 9.465 0.405 ;
        RECT  8.575 -0.250 9.205 0.250 ;
        RECT  8.315 -0.250 8.575 0.405 ;
        RECT  7.135 -0.250 8.315 0.250 ;
        RECT  6.875 -0.250 7.135 0.405 ;
        RECT  5.580 -0.250 6.875 0.250 ;
        RECT  5.320 -0.250 5.580 0.405 ;
        RECT  4.715 -0.250 5.320 0.250 ;
        RECT  4.455 -0.250 4.715 0.405 ;
        RECT  3.440 -0.250 4.455 0.250 ;
        RECT  3.180 -0.250 3.440 0.405 ;
        RECT  0.815 -0.250 3.180 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.620 3.440 14.720 3.940 ;
        RECT  13.360 2.610 13.620 3.940 ;
        RECT  11.645 3.440 13.360 3.940 ;
        RECT  11.385 3.285 11.645 3.940 ;
        RECT  6.945 3.440 11.385 3.940 ;
        RECT  6.685 3.285 6.945 3.940 ;
        RECT  4.825 3.440 6.685 3.940 ;
        RECT  4.565 2.945 4.825 3.940 ;
        RECT  3.815 3.440 4.565 3.940 ;
        RECT  3.555 2.945 3.815 3.940 ;
        RECT  2.575 3.440 3.555 3.940 ;
        RECT  2.315 2.780 2.575 3.940 ;
        RECT  0.815 3.440 2.315 3.940 ;
        RECT  0.555 3.285 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.055 2.000 14.200 2.260 ;
        RECT  14.055 0.430 14.175 0.590 ;
        RECT  14.040 0.430 14.055 2.260 ;
        RECT  13.895 0.430 14.040 2.160 ;
        RECT  12.785 0.585 13.895 0.745 ;
        RECT  13.400 2.000 13.895 2.160 ;
        RECT  13.550 1.380 13.710 1.645 ;
        RECT  13.370 1.380 13.550 1.540 ;
        RECT  13.240 1.895 13.400 2.160 ;
        RECT  13.210 0.925 13.370 1.540 ;
        RECT  12.535 0.925 13.210 1.085 ;
        RECT  12.995 2.975 13.080 3.235 ;
        RECT  12.835 1.265 12.995 3.235 ;
        RECT  12.760 1.265 12.835 1.525 ;
        RECT  12.820 2.915 12.835 3.235 ;
        RECT  10.855 2.915 12.820 3.075 ;
        RECT  12.625 0.470 12.785 0.745 ;
        RECT  12.535 2.410 12.655 2.670 ;
        RECT  9.805 0.470 12.625 0.630 ;
        RECT  12.375 0.925 12.535 2.670 ;
        RECT  12.360 1.130 12.375 1.390 ;
        RECT  12.090 2.475 12.195 2.735 ;
        RECT  10.150 0.810 12.180 0.970 ;
        RECT  11.930 1.195 12.090 2.735 ;
        RECT  11.660 1.195 11.930 1.355 ;
        RECT  11.165 2.575 11.930 2.735 ;
        RECT  11.235 1.845 11.750 2.105 ;
        RECT  11.075 1.185 11.235 2.395 ;
        RECT  10.330 1.185 11.075 1.345 ;
        RECT  10.695 2.235 11.075 2.395 ;
        RECT  10.355 1.890 10.895 2.050 ;
        RECT  10.695 2.720 10.855 3.075 ;
        RECT  10.535 2.235 10.695 2.540 ;
        RECT  10.355 2.720 10.695 2.880 ;
        RECT  7.285 3.060 10.515 3.220 ;
        RECT  10.195 1.545 10.355 2.880 ;
        RECT  9.760 1.545 10.195 1.705 ;
        RECT  7.625 2.720 10.195 2.880 ;
        RECT  9.990 0.810 10.150 1.150 ;
        RECT  9.390 1.895 10.015 2.055 ;
        RECT  9.390 0.990 9.990 1.150 ;
        RECT  9.645 0.470 9.805 0.760 ;
        RECT  9.600 1.365 9.760 1.705 ;
        RECT  6.875 0.600 9.645 0.760 ;
        RECT  9.230 0.990 9.390 2.540 ;
        RECT  8.850 0.990 9.230 1.250 ;
        RECT  7.965 2.380 9.230 2.540 ;
        RECT  8.420 1.500 9.050 1.760 ;
        RECT  8.260 1.135 8.420 2.165 ;
        RECT  8.140 1.135 8.260 1.295 ;
        RECT  8.160 2.005 8.260 2.165 ;
        RECT  7.880 1.035 8.140 1.295 ;
        RECT  7.805 2.125 7.965 2.540 ;
        RECT  7.465 2.605 7.625 2.880 ;
        RECT  7.265 0.950 7.610 1.110 ;
        RECT  7.265 2.605 7.465 2.765 ;
        RECT  7.125 2.945 7.285 3.220 ;
        RECT  7.105 0.950 7.265 2.765 ;
        RECT  6.505 2.945 7.125 3.105 ;
        RECT  6.715 0.600 6.875 1.720 ;
        RECT  6.505 2.150 6.535 2.410 ;
        RECT  6.345 0.720 6.505 3.220 ;
        RECT  6.245 0.720 6.345 0.880 ;
        RECT  5.165 3.060 6.345 3.220 ;
        RECT  5.985 0.620 6.245 0.880 ;
        RECT  6.005 1.180 6.165 2.875 ;
        RECT  5.900 1.180 6.005 1.340 ;
        RECT  5.735 2.715 6.005 2.875 ;
        RECT  5.655 1.500 5.795 1.760 ;
        RECT  5.495 1.085 5.655 2.295 ;
        RECT  4.890 1.085 5.495 1.245 ;
        RECT  5.275 2.135 5.495 2.295 ;
        RECT  5.005 2.605 5.165 3.220 ;
        RECT  2.915 2.605 5.005 2.765 ;
        RECT  3.605 2.240 4.245 2.400 ;
        RECT  3.605 1.085 3.815 1.245 ;
        RECT  3.445 1.085 3.605 2.400 ;
        RECT  3.155 1.590 3.445 1.850 ;
        RECT  2.975 1.130 3.255 1.390 ;
        RECT  2.975 2.100 3.255 2.260 ;
        RECT  2.815 1.130 2.975 2.260 ;
        RECT  2.755 2.440 2.915 2.765 ;
        RECT  2.635 1.130 2.815 1.290 ;
        RECT  1.655 2.440 2.755 2.600 ;
        RECT  2.475 0.810 2.635 1.290 ;
        RECT  1.835 0.810 2.475 0.970 ;
        RECT  2.115 1.180 2.295 1.340 ;
        RECT  2.115 2.100 2.215 2.260 ;
        RECT  1.955 1.180 2.115 2.260 ;
        RECT  1.505 2.780 1.765 3.035 ;
        RECT  1.495 1.130 1.655 2.600 ;
        RECT  0.385 2.780 1.505 2.940 ;
        RECT  0.325 2.255 0.385 2.940 ;
        RECT  0.325 1.025 0.335 1.285 ;
        RECT  0.225 1.025 0.325 2.940 ;
        RECT  0.165 1.025 0.225 2.515 ;
        RECT  0.125 2.255 0.165 2.515 ;
    END
END SEDFFHQX1

MACRO SDFFSRHQX8
    CLASS CORE ;
    FOREIGN SDFFSRHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.320 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.655 7.695 2.400 ;
        RECT  7.435 1.655 7.485 1.915 ;
        END
        ANTENNAGATEAREA     0.2691 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.185 1.265 6.375 2.080 ;
        RECT  5.965 1.265 6.185 1.635 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.340 1.615 5.445 1.875 ;
        RECT  5.180 1.615 5.340 2.540 ;
        RECT  2.755 2.380 5.180 2.540 ;
        RECT  2.595 1.620 2.755 2.540 ;
        RECT  2.425 1.700 2.595 2.175 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.165 1.525 14.425 1.785 ;
        RECT  13.215 1.625 14.165 1.785 ;
        RECT  12.845 1.625 13.215 1.990 ;
        END
        ANTENNAGATEAREA     0.3419 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.735 0.980 19.195 2.395 ;
        RECT  18.685 0.980 18.735 2.585 ;
        RECT  18.525 0.690 18.685 3.045 ;
        RECT  18.425 0.690 18.525 1.290 ;
        RECT  18.425 1.990 18.525 3.045 ;
        RECT  17.665 0.980 18.425 1.290 ;
        RECT  18.275 1.990 18.425 2.400 ;
        RECT  17.665 1.990 18.275 2.395 ;
        RECT  17.405 0.690 17.665 1.290 ;
        RECT  17.405 1.990 17.665 3.045 ;
        END
        ANTENNADIFFAREA     1.6264 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.625 1.290 4.265 1.580 ;
        END
        ANTENNAGATEAREA     0.2366 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.335 2.185 ;
        END
        ANTENNAGATEAREA     0.3783 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.195 -0.250 19.320 0.250 ;
        RECT  18.935 -0.250 19.195 0.755 ;
        RECT  18.175 -0.250 18.935 0.250 ;
        RECT  17.915 -0.250 18.175 0.755 ;
        RECT  17.125 -0.250 17.915 0.250 ;
        RECT  16.865 -0.250 17.125 1.135 ;
        RECT  16.525 -0.250 16.865 0.405 ;
        RECT  15.115 -0.250 16.525 0.250 ;
        RECT  14.855 -0.250 15.115 0.405 ;
        RECT  12.070 -0.250 14.855 0.250 ;
        RECT  11.810 -0.250 12.070 0.405 ;
        RECT  9.830 -0.250 11.810 0.250 ;
        RECT  9.230 -0.250 9.830 0.405 ;
        RECT  7.615 -0.250 9.230 0.250 ;
        RECT  7.355 -0.250 7.615 0.405 ;
        RECT  6.595 -0.250 7.355 0.250 ;
        RECT  5.995 -0.250 6.595 0.405 ;
        RECT  4.115 -0.250 5.995 0.250 ;
        RECT  3.875 -0.250 4.115 0.405 ;
        RECT  3.515 -0.250 3.875 0.745 ;
        RECT  0.940 -0.250 3.515 0.250 ;
        RECT  0.340 -0.250 0.940 0.405 ;
        RECT  0.000 -0.250 0.340 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.195 3.440 19.320 3.940 ;
        RECT  18.935 2.615 19.195 3.940 ;
        RECT  18.175 3.440 18.935 3.940 ;
        RECT  17.915 2.615 18.175 3.940 ;
        RECT  17.155 3.440 17.915 3.940 ;
        RECT  16.895 2.275 17.155 3.940 ;
        RECT  16.215 2.955 16.895 3.940 ;
        RECT  14.775 3.440 16.215 3.940 ;
        RECT  14.515 3.285 14.775 3.940 ;
        RECT  12.135 3.440 14.515 3.940 ;
        RECT  11.875 3.285 12.135 3.940 ;
        RECT  10.990 3.440 11.875 3.940 ;
        RECT  10.730 3.285 10.990 3.940 ;
        RECT  9.460 3.440 10.730 3.940 ;
        RECT  9.200 2.660 9.460 3.940 ;
        RECT  6.920 3.440 9.200 3.940 ;
        RECT  6.660 3.285 6.920 3.940 ;
        RECT  1.380 3.440 6.660 3.940 ;
        RECT  0.780 3.285 1.380 3.940 ;
        RECT  0.000 3.440 0.780 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.325 1.510 18.055 1.770 ;
        RECT  16.665 1.495 17.325 1.770 ;
        RECT  16.505 0.680 16.665 2.580 ;
        RECT  15.655 0.680 16.505 0.840 ;
        RECT  16.435 1.510 16.505 1.770 ;
        RECT  15.725 2.420 16.505 2.580 ;
        RECT  16.225 1.035 16.325 1.295 ;
        RECT  16.225 1.955 16.325 2.215 ;
        RECT  16.065 1.035 16.225 2.215 ;
        RECT  15.695 1.725 16.065 1.985 ;
        RECT  15.565 2.420 15.725 2.935 ;
        RECT  15.495 0.680 15.655 1.025 ;
        RECT  13.825 2.775 15.565 2.935 ;
        RECT  15.395 0.765 15.495 1.025 ;
        RECT  15.385 1.205 15.485 1.465 ;
        RECT  13.315 0.840 15.395 1.000 ;
        RECT  15.285 1.205 15.385 2.295 ;
        RECT  15.225 1.205 15.285 2.595 ;
        RECT  15.125 2.035 15.225 2.595 ;
        RECT  14.115 2.435 15.125 2.595 ;
        RECT  14.805 1.995 14.905 2.255 ;
        RECT  14.645 1.180 14.805 2.255 ;
        RECT  13.095 1.180 14.645 1.340 ;
        RECT  13.955 2.055 14.115 2.595 ;
        RECT  13.825 2.055 13.955 2.330 ;
        RECT  13.095 0.470 13.945 0.630 ;
        RECT  12.665 2.170 13.825 2.330 ;
        RECT  13.565 2.775 13.825 3.035 ;
        RECT  12.660 2.510 13.260 2.770 ;
        RECT  12.935 0.470 13.095 1.340 ;
        RECT  12.475 3.060 13.055 3.220 ;
        RECT  12.415 0.470 12.935 0.630 ;
        RECT  12.665 0.810 12.755 1.085 ;
        RECT  12.595 0.810 12.665 2.330 ;
        RECT  11.585 2.510 12.660 2.670 ;
        RECT  12.505 0.925 12.595 2.330 ;
        RECT  11.290 0.925 12.505 1.085 ;
        RECT  12.005 2.015 12.505 2.330 ;
        RECT  12.315 2.945 12.475 3.220 ;
        RECT  12.255 0.470 12.415 0.745 ;
        RECT  12.155 1.265 12.315 1.525 ;
        RECT  10.450 2.945 12.315 3.105 ;
        RECT  11.630 0.585 12.255 0.745 ;
        RECT  10.950 1.265 12.155 1.425 ;
        RECT  11.470 0.470 11.630 0.745 ;
        RECT  11.325 2.460 11.585 2.720 ;
        RECT  10.170 0.470 11.470 0.630 ;
        RECT  10.960 2.460 11.325 2.620 ;
        RECT  11.130 0.810 11.290 1.085 ;
        RECT  10.510 0.810 11.130 0.970 ;
        RECT  10.950 1.920 10.960 2.620 ;
        RECT  10.800 1.150 10.950 2.620 ;
        RECT  10.790 1.150 10.800 2.130 ;
        RECT  10.690 1.150 10.790 1.425 ;
        RECT  10.675 1.870 10.790 2.130 ;
        RECT  10.350 0.810 10.510 1.145 ;
        RECT  10.350 1.385 10.510 1.645 ;
        RECT  10.190 2.945 10.450 3.245 ;
        RECT  7.250 0.985 10.350 1.145 ;
        RECT  10.230 1.485 10.350 1.645 ;
        RECT  10.230 2.390 10.280 2.650 ;
        RECT  10.070 1.485 10.230 2.650 ;
        RECT  9.800 2.945 10.190 3.105 ;
        RECT  10.010 0.470 10.170 0.745 ;
        RECT  9.075 1.485 10.070 1.645 ;
        RECT  10.020 2.390 10.070 2.650 ;
        RECT  9.335 0.585 10.010 0.745 ;
        RECT  9.640 2.210 9.800 3.105 ;
        RECT  8.720 2.210 9.640 2.370 ;
        RECT  9.075 0.585 9.335 0.805 ;
        RECT  4.215 0.585 9.075 0.745 ;
        RECT  8.815 1.325 9.075 1.645 ;
        RECT  8.035 1.485 8.815 1.645 ;
        RECT  8.560 1.925 8.720 3.220 ;
        RECT  8.375 1.925 8.560 2.085 ;
        RECT  7.260 3.060 8.560 3.220 ;
        RECT  7.600 2.720 8.380 2.880 ;
        RECT  8.215 1.825 8.375 2.085 ;
        RECT  8.035 2.350 8.240 2.510 ;
        RECT  7.875 1.485 8.035 2.510 ;
        RECT  7.440 2.605 7.600 2.880 ;
        RECT  6.715 2.605 7.440 2.765 ;
        RECT  7.250 2.265 7.290 2.425 ;
        RECT  7.100 2.945 7.260 3.220 ;
        RECT  7.090 0.935 7.250 2.425 ;
        RECT  6.480 2.945 7.100 3.105 ;
        RECT  6.895 0.935 7.090 1.195 ;
        RECT  7.030 2.265 7.090 2.425 ;
        RECT  6.555 0.925 6.715 2.765 ;
        RECT  5.215 0.925 6.555 1.085 ;
        RECT  5.860 2.395 6.555 2.655 ;
        RECT  6.320 2.945 6.480 3.220 ;
        RECT  1.725 3.060 6.320 3.220 ;
        RECT  5.785 1.865 6.005 2.215 ;
        RECT  5.680 1.275 5.785 2.215 ;
        RECT  5.625 1.275 5.680 2.880 ;
        RECT  4.965 1.275 5.625 1.435 ;
        RECT  5.520 2.055 5.625 2.880 ;
        RECT  2.235 2.720 5.520 2.880 ;
        RECT  4.955 0.925 5.215 1.095 ;
        RECT  4.605 2.040 5.000 2.200 ;
        RECT  4.785 1.275 4.965 1.560 ;
        RECT  4.605 0.925 4.655 1.085 ;
        RECT  4.445 0.925 4.605 2.200 ;
        RECT  4.395 0.925 4.445 1.085 ;
        RECT  4.055 0.585 4.215 1.110 ;
        RECT  3.235 0.950 4.055 1.110 ;
        RECT  3.235 2.040 4.050 2.200 ;
        RECT  3.075 0.930 3.235 2.200 ;
        RECT  2.975 0.930 3.075 1.190 ;
        RECT  2.765 0.470 2.975 0.750 ;
        RECT  2.575 0.930 2.975 1.090 ;
        RECT  1.285 0.470 2.765 0.630 ;
        RECT  2.415 0.810 2.575 1.090 ;
        RECT  1.625 0.810 2.415 0.970 ;
        RECT  2.075 1.150 2.235 2.880 ;
        RECT  1.805 1.150 2.075 1.310 ;
        RECT  1.625 1.575 1.895 1.835 ;
        RECT  1.565 2.120 1.725 3.220 ;
        RECT  1.465 0.810 1.625 1.835 ;
        RECT  1.465 2.120 1.565 2.380 ;
        RECT  1.295 1.575 1.465 1.835 ;
        RECT  1.015 2.120 1.465 2.280 ;
        RECT  1.125 0.470 1.285 0.745 ;
        RECT  1.125 0.970 1.285 1.230 ;
        RECT  0.675 0.585 1.125 0.745 ;
        RECT  1.015 1.070 1.125 1.230 ;
        RECT  0.855 1.070 1.015 2.280 ;
        RECT  0.515 0.585 0.675 2.895 ;
        RECT  0.125 0.835 0.515 1.095 ;
        RECT  0.385 2.735 0.515 2.895 ;
        RECT  0.125 2.735 0.385 2.995 ;
    END
END SDFFSRHQX8

MACRO SDFFSRHQX4
    CLASS CORE ;
    FOREIGN SDFFSRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.940 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.655 7.695 2.400 ;
        RECT  7.435 1.655 7.485 1.915 ;
        END
        ANTENNAGATEAREA     0.2691 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.185 1.265 6.375 2.080 ;
        RECT  5.965 1.265 6.185 1.635 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.340 1.615 5.445 1.875 ;
        RECT  5.180 1.615 5.340 2.540 ;
        RECT  2.755 2.380 5.180 2.540 ;
        RECT  2.595 1.620 2.755 2.540 ;
        RECT  2.425 1.700 2.595 2.175 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.295 1.525 14.455 1.820 ;
        RECT  13.215 1.660 14.295 1.820 ;
        RECT  13.125 1.660 13.215 1.990 ;
        RECT  13.005 1.585 13.125 1.990 ;
        RECT  12.965 1.585 13.005 1.845 ;
        END
        ANTENNAGATEAREA     0.3419 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.605 1.080 17.815 2.315 ;
        RECT  17.295 1.080 17.605 1.290 ;
        RECT  17.355 2.105 17.605 2.315 ;
        RECT  17.295 2.105 17.355 2.585 ;
        RECT  17.035 0.690 17.295 1.290 ;
        RECT  17.035 2.105 17.295 3.045 ;
        END
        ANTENNADIFFAREA     0.8132 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.625 1.290 4.265 1.580 ;
        END
        ANTENNAGATEAREA     0.2366 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.335 2.185 ;
        END
        ANTENNAGATEAREA     0.3783 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.805 -0.250 17.940 0.250 ;
        RECT  17.545 -0.250 17.805 0.755 ;
        RECT  16.755 -0.250 17.545 0.250 ;
        RECT  16.495 -0.250 16.755 0.405 ;
        RECT  15.195 -0.250 16.495 0.250 ;
        RECT  14.935 -0.250 15.195 0.405 ;
        RECT  12.070 -0.250 14.935 0.250 ;
        RECT  11.810 -0.250 12.070 0.405 ;
        RECT  9.830 -0.250 11.810 0.250 ;
        RECT  9.230 -0.250 9.830 0.405 ;
        RECT  7.615 -0.250 9.230 0.250 ;
        RECT  7.355 -0.250 7.615 0.405 ;
        RECT  6.595 -0.250 7.355 0.250 ;
        RECT  5.995 -0.250 6.595 0.405 ;
        RECT  4.115 -0.250 5.995 0.250 ;
        RECT  3.875 -0.250 4.115 0.405 ;
        RECT  3.515 -0.250 3.875 0.745 ;
        RECT  0.940 -0.250 3.515 0.250 ;
        RECT  0.340 -0.250 0.940 0.405 ;
        RECT  0.000 -0.250 0.340 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.805 3.440 17.940 3.940 ;
        RECT  17.545 2.615 17.805 3.940 ;
        RECT  16.785 3.440 17.545 3.940 ;
        RECT  16.185 2.955 16.785 3.940 ;
        RECT  14.775 3.440 16.185 3.940 ;
        RECT  14.515 3.285 14.775 3.940 ;
        RECT  12.135 3.440 14.515 3.940 ;
        RECT  11.875 3.285 12.135 3.940 ;
        RECT  10.990 3.440 11.875 3.940 ;
        RECT  10.730 3.285 10.990 3.940 ;
        RECT  9.460 3.440 10.730 3.940 ;
        RECT  9.200 2.660 9.460 3.940 ;
        RECT  6.920 3.440 9.200 3.940 ;
        RECT  6.660 3.285 6.920 3.940 ;
        RECT  1.380 3.440 6.660 3.940 ;
        RECT  0.780 3.285 1.380 3.940 ;
        RECT  0.000 3.440 0.780 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.695 1.495 17.375 1.755 ;
        RECT  16.665 0.695 16.695 1.755 ;
        RECT  16.535 0.695 16.665 2.580 ;
        RECT  15.735 0.695 16.535 0.855 ;
        RECT  16.505 1.495 16.535 2.580 ;
        RECT  16.435 1.495 16.505 1.755 ;
        RECT  15.725 2.420 16.505 2.580 ;
        RECT  16.225 1.035 16.325 1.295 ;
        RECT  16.225 1.955 16.325 2.215 ;
        RECT  16.065 1.035 16.225 2.215 ;
        RECT  15.605 1.725 16.065 1.985 ;
        RECT  15.475 0.695 15.735 1.035 ;
        RECT  15.565 2.420 15.725 2.935 ;
        RECT  13.825 2.775 15.565 2.935 ;
        RECT  13.565 0.840 15.475 1.000 ;
        RECT  15.385 1.215 15.415 1.475 ;
        RECT  15.285 1.215 15.385 2.295 ;
        RECT  15.225 1.215 15.285 2.595 ;
        RECT  15.155 1.215 15.225 1.475 ;
        RECT  15.125 2.035 15.225 2.595 ;
        RECT  14.085 2.435 15.125 2.595 ;
        RECT  14.750 1.180 14.910 2.215 ;
        RECT  13.350 1.180 14.750 1.340 ;
        RECT  14.645 2.055 14.750 2.215 ;
        RECT  13.350 0.470 14.085 0.630 ;
        RECT  13.925 2.005 14.085 2.595 ;
        RECT  13.825 2.005 13.925 2.330 ;
        RECT  12.750 2.170 13.825 2.330 ;
        RECT  13.565 2.775 13.825 3.035 ;
        RECT  13.190 0.470 13.350 1.340 ;
        RECT  12.660 2.515 13.260 2.775 ;
        RECT  12.410 0.470 13.190 0.630 ;
        RECT  12.475 3.060 13.055 3.220 ;
        RECT  12.750 0.810 12.850 1.070 ;
        RECT  12.590 0.810 12.750 2.330 ;
        RECT  10.950 2.605 12.660 2.765 ;
        RECT  11.290 0.925 12.590 1.085 ;
        RECT  12.265 2.065 12.590 2.225 ;
        RECT  12.315 2.945 12.475 3.220 ;
        RECT  12.250 0.470 12.410 0.745 ;
        RECT  10.950 1.265 12.405 1.425 ;
        RECT  10.450 2.945 12.315 3.105 ;
        RECT  12.005 2.015 12.265 2.275 ;
        RECT  11.630 0.585 12.250 0.745 ;
        RECT  11.470 0.470 11.630 0.745 ;
        RECT  10.170 0.470 11.470 0.630 ;
        RECT  11.130 0.810 11.290 1.085 ;
        RECT  10.510 0.810 11.130 0.970 ;
        RECT  10.790 1.150 10.950 2.765 ;
        RECT  10.690 1.150 10.790 1.425 ;
        RECT  10.675 1.870 10.790 2.130 ;
        RECT  10.350 0.810 10.510 1.145 ;
        RECT  10.350 1.385 10.510 1.645 ;
        RECT  10.190 2.945 10.450 3.260 ;
        RECT  7.250 0.985 10.350 1.145 ;
        RECT  10.230 1.485 10.350 1.645 ;
        RECT  10.230 2.605 10.280 2.765 ;
        RECT  10.070 1.485 10.230 2.765 ;
        RECT  9.800 2.945 10.190 3.105 ;
        RECT  10.010 0.470 10.170 0.745 ;
        RECT  9.075 1.485 10.070 1.645 ;
        RECT  10.020 2.605 10.070 2.765 ;
        RECT  9.335 0.585 10.010 0.745 ;
        RECT  9.640 2.210 9.800 3.105 ;
        RECT  8.720 2.210 9.640 2.370 ;
        RECT  9.075 0.585 9.335 0.805 ;
        RECT  4.215 0.585 9.075 0.745 ;
        RECT  8.815 1.325 9.075 1.645 ;
        RECT  8.035 1.485 8.815 1.645 ;
        RECT  8.560 1.925 8.720 3.220 ;
        RECT  8.375 1.925 8.560 2.085 ;
        RECT  7.260 3.060 8.560 3.220 ;
        RECT  7.600 2.720 8.380 2.880 ;
        RECT  8.215 1.825 8.375 2.085 ;
        RECT  8.035 2.350 8.240 2.510 ;
        RECT  7.875 1.485 8.035 2.510 ;
        RECT  7.440 2.605 7.600 2.880 ;
        RECT  6.715 2.605 7.440 2.765 ;
        RECT  7.250 2.265 7.290 2.425 ;
        RECT  7.100 2.945 7.260 3.220 ;
        RECT  7.090 0.935 7.250 2.425 ;
        RECT  6.480 2.945 7.100 3.105 ;
        RECT  6.895 0.935 7.090 1.195 ;
        RECT  7.030 2.265 7.090 2.425 ;
        RECT  6.555 0.925 6.715 2.765 ;
        RECT  5.215 0.925 6.555 1.085 ;
        RECT  5.860 2.395 6.555 2.655 ;
        RECT  6.320 2.945 6.480 3.220 ;
        RECT  1.725 3.060 6.320 3.220 ;
        RECT  5.785 1.865 6.005 2.215 ;
        RECT  5.680 1.275 5.785 2.215 ;
        RECT  5.625 1.275 5.680 2.880 ;
        RECT  4.965 1.275 5.625 1.435 ;
        RECT  5.520 2.055 5.625 2.880 ;
        RECT  2.235 2.720 5.520 2.880 ;
        RECT  4.955 0.925 5.215 1.095 ;
        RECT  4.605 2.040 5.000 2.200 ;
        RECT  4.785 1.275 4.965 1.560 ;
        RECT  4.605 0.925 4.655 1.085 ;
        RECT  4.445 0.925 4.605 2.200 ;
        RECT  4.395 0.925 4.445 1.085 ;
        RECT  4.055 0.585 4.215 1.110 ;
        RECT  3.235 0.950 4.055 1.110 ;
        RECT  3.235 2.040 4.050 2.200 ;
        RECT  3.075 0.930 3.235 2.200 ;
        RECT  2.975 0.930 3.075 1.190 ;
        RECT  2.765 0.470 2.975 0.750 ;
        RECT  2.575 0.930 2.975 1.090 ;
        RECT  1.285 0.470 2.765 0.630 ;
        RECT  2.415 0.810 2.575 1.090 ;
        RECT  1.625 0.810 2.415 0.970 ;
        RECT  2.075 1.150 2.235 2.880 ;
        RECT  1.805 1.150 2.075 1.310 ;
        RECT  1.625 1.575 1.895 1.835 ;
        RECT  1.565 2.120 1.725 3.220 ;
        RECT  1.465 0.810 1.625 1.835 ;
        RECT  1.465 2.120 1.565 2.380 ;
        RECT  1.295 1.575 1.465 1.835 ;
        RECT  1.015 2.120 1.465 2.280 ;
        RECT  1.125 0.470 1.285 0.745 ;
        RECT  1.125 0.970 1.285 1.230 ;
        RECT  0.675 0.585 1.125 0.745 ;
        RECT  1.015 1.070 1.125 1.230 ;
        RECT  0.855 1.070 1.015 2.280 ;
        RECT  0.515 0.585 0.675 2.895 ;
        RECT  0.125 0.835 0.515 1.095 ;
        RECT  0.385 2.735 0.515 2.895 ;
        RECT  0.125 2.735 0.385 2.995 ;
    END
END SDFFSRHQX4

MACRO SDFFSRHQX2
    CLASS CORE ;
    FOREIGN SDFFSRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.100 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.285 1.580 6.775 1.990 ;
        END
        ANTENNAGATEAREA     0.1911 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.035 1.290 5.395 1.845 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.355 1.805 4.515 2.425 ;
        RECT  2.635 2.265 4.355 2.425 ;
        RECT  2.425 2.110 2.635 2.425 ;
        RECT  2.315 2.165 2.425 2.425 ;
        END
        ANTENNAGATEAREA     0.1833 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.755 1.665 12.830 1.925 ;
        RECT  12.570 1.665 12.755 1.990 ;
        RECT  12.545 1.700 12.570 1.990 ;
        RECT  11.955 1.715 12.545 1.875 ;
        RECT  11.795 1.715 11.955 2.055 ;
        RECT  10.795 1.895 11.795 2.055 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.715 0.695 15.975 1.450 ;
        RECT  15.515 1.290 15.715 1.450 ;
        RECT  15.515 1.925 15.545 2.555 ;
        RECT  15.305 1.290 15.515 2.555 ;
        RECT  15.285 1.955 15.305 2.555 ;
        END
        ANTENNADIFFAREA     0.5668 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.225 1.155 3.635 1.580 ;
        END
        ANTENNAGATEAREA     0.1677 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.795 1.845 ;
        RECT  0.535 1.585 0.585 1.845 ;
        END
        ANTENNAGATEAREA     0.2314 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.435 -0.250 16.100 0.250 ;
        RECT  15.175 -0.250 15.435 1.090 ;
        RECT  14.835 -0.250 15.175 0.405 ;
        RECT  13.520 -0.250 14.835 0.250 ;
        RECT  13.260 -0.250 13.520 0.405 ;
        RECT  9.065 -0.250 13.260 0.250 ;
        RECT  8.805 -0.250 9.065 0.405 ;
        RECT  5.975 -0.250 8.805 0.250 ;
        RECT  5.715 -0.250 5.975 0.405 ;
        RECT  3.145 -0.250 5.715 0.250 ;
        RECT  2.885 -0.250 3.145 0.405 ;
        RECT  0.935 -0.250 2.885 0.250 ;
        RECT  0.675 -0.250 0.935 0.405 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.945 3.440 16.100 3.940 ;
        RECT  14.885 3.285 15.945 3.940 ;
        RECT  12.935 3.440 14.885 3.940 ;
        RECT  12.675 3.285 12.935 3.940 ;
        RECT  10.515 3.440 12.675 3.940 ;
        RECT  10.255 3.285 10.515 3.940 ;
        RECT  9.565 3.440 10.255 3.940 ;
        RECT  9.305 3.285 9.565 3.940 ;
        RECT  8.315 3.440 9.305 3.940 ;
        RECT  8.055 3.285 8.315 3.940 ;
        RECT  6.005 3.440 8.055 3.940 ;
        RECT  5.745 3.285 6.005 3.940 ;
        RECT  3.775 3.440 5.745 3.940 ;
        RECT  3.515 3.285 3.775 3.940 ;
        RECT  1.405 3.440 3.515 3.940 ;
        RECT  0.725 3.285 1.405 3.940 ;
        RECT  0.465 2.890 0.725 3.940 ;
        RECT  0.000 3.440 0.465 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.975 1.580 15.105 1.840 ;
        RECT  14.815 0.675 14.975 3.085 ;
        RECT  14.095 0.675 14.815 0.835 ;
        RECT  12.200 2.925 14.815 3.085 ;
        RECT  14.425 2.465 14.635 2.725 ;
        RECT  14.425 1.035 14.525 1.295 ;
        RECT  14.265 1.035 14.425 2.725 ;
        RECT  14.005 1.495 14.265 1.755 ;
        RECT  13.835 0.525 14.095 0.835 ;
        RECT  13.785 1.015 14.005 1.275 ;
        RECT  12.320 0.675 13.835 0.835 ;
        RECT  13.685 1.015 13.785 2.450 ;
        RECT  13.625 1.015 13.685 2.745 ;
        RECT  13.525 2.190 13.625 2.745 ;
        RECT  12.540 2.585 13.525 2.745 ;
        RECT  13.255 2.145 13.305 2.405 ;
        RECT  13.095 1.235 13.255 2.405 ;
        RECT  11.880 1.235 13.095 1.395 ;
        RECT  13.045 2.145 13.095 2.405 ;
        RECT  12.395 2.265 12.540 2.745 ;
        RECT  12.380 2.165 12.395 2.745 ;
        RECT  12.135 2.165 12.380 2.425 ;
        RECT  12.060 0.675 12.320 1.055 ;
        RECT  12.040 2.655 12.200 3.085 ;
        RECT  10.610 2.265 12.135 2.425 ;
        RECT  11.940 2.655 12.040 2.915 ;
        RECT  11.720 0.470 11.880 1.395 ;
        RECT  9.405 0.470 11.720 0.630 ;
        RECT  11.205 2.605 11.465 2.885 ;
        RECT  11.255 0.810 11.415 1.715 ;
        RECT  11.025 3.065 11.365 3.225 ;
        RECT  9.745 0.810 11.255 0.970 ;
        RECT  10.610 1.555 11.255 1.715 ;
        RECT  10.115 2.605 11.205 2.765 ;
        RECT  10.130 1.205 11.075 1.365 ;
        RECT  10.865 2.945 11.025 3.225 ;
        RECT  9.025 2.945 10.865 3.105 ;
        RECT  10.450 1.555 10.610 2.425 ;
        RECT  10.315 2.265 10.450 2.425 ;
        RECT  9.970 1.205 10.130 1.425 ;
        RECT  9.955 2.185 10.115 2.765 ;
        RECT  9.470 1.265 9.970 1.425 ;
        RECT  9.470 2.185 9.955 2.345 ;
        RECT  9.585 0.810 9.745 1.085 ;
        RECT  8.285 0.925 9.585 1.085 ;
        RECT  9.310 1.265 9.470 2.345 ;
        RECT  9.245 0.470 9.405 0.745 ;
        RECT  9.075 1.935 9.310 2.195 ;
        RECT  8.625 0.585 9.245 0.745 ;
        RECT  8.895 1.455 9.130 1.715 ;
        RECT  8.765 2.945 9.025 3.205 ;
        RECT  8.735 1.455 8.895 2.760 ;
        RECT  7.235 2.945 8.765 3.105 ;
        RECT  8.565 2.500 8.735 2.760 ;
        RECT  8.465 0.470 8.625 0.745 ;
        RECT  7.555 2.600 8.565 2.760 ;
        RECT  6.315 0.470 8.465 0.630 ;
        RECT  8.125 0.810 8.285 1.085 ;
        RECT  6.655 0.810 8.125 0.970 ;
        RECT  7.765 1.150 7.945 1.310 ;
        RECT  7.605 1.150 7.765 2.270 ;
        RECT  7.555 2.110 7.605 2.270 ;
        RECT  7.395 2.110 7.555 2.760 ;
        RECT  7.215 1.445 7.265 1.705 ;
        RECT  7.215 2.945 7.235 3.210 ;
        RECT  7.055 1.445 7.215 3.210 ;
        RECT  7.005 1.445 7.055 1.705 ;
        RECT  6.345 3.050 7.055 3.210 ;
        RECT  6.715 2.555 6.875 2.870 ;
        RECT  5.735 2.555 6.715 2.715 ;
        RECT  6.495 0.810 6.655 1.110 ;
        RECT  6.075 0.950 6.495 1.110 ;
        RECT  6.185 2.945 6.345 3.210 ;
        RECT  6.155 0.470 6.315 0.745 ;
        RECT  3.045 2.945 6.185 3.105 ;
        RECT  5.535 0.585 6.155 0.745 ;
        RECT  5.915 0.950 6.075 2.255 ;
        RECT  5.575 0.925 5.735 2.715 ;
        RECT  5.195 0.925 5.575 1.085 ;
        RECT  5.195 2.505 5.575 2.715 ;
        RECT  5.375 0.475 5.535 0.745 ;
        RECT  4.855 2.115 5.390 2.275 ;
        RECT  3.485 0.475 5.375 0.635 ;
        RECT  5.035 0.815 5.195 1.085 ;
        RECT  5.035 2.505 5.195 2.765 ;
        RECT  4.225 0.815 5.035 0.975 ;
        RECT  4.695 1.335 4.855 2.765 ;
        RECT  4.315 1.335 4.695 1.495 ;
        RECT  2.705 2.605 4.695 2.765 ;
        RECT  4.155 1.155 4.315 1.495 ;
        RECT  3.975 1.925 4.175 2.085 ;
        RECT  3.815 0.815 3.975 2.085 ;
        RECT  3.715 0.815 3.815 0.975 ;
        RECT  3.325 0.475 3.485 0.970 ;
        RECT  2.975 0.810 3.325 0.970 ;
        RECT  2.975 1.925 3.225 2.085 ;
        RECT  2.885 2.945 3.045 3.220 ;
        RECT  2.815 0.810 2.975 2.085 ;
        RECT  1.765 3.060 2.885 3.220 ;
        RECT  2.555 0.810 2.815 1.075 ;
        RECT  2.445 2.605 2.705 2.880 ;
        RECT  1.705 0.810 2.555 0.970 ;
        RECT  2.135 2.605 2.445 2.765 ;
        RECT  2.135 1.150 2.305 1.310 ;
        RECT  1.310 0.460 2.145 0.620 ;
        RECT  1.975 1.150 2.135 2.765 ;
        RECT  1.605 2.070 1.765 3.220 ;
        RECT  1.545 0.810 1.705 1.845 ;
        RECT  1.505 2.070 1.605 2.670 ;
        RECT  1.335 1.585 1.545 1.845 ;
        RECT  1.135 2.070 1.505 2.230 ;
        RECT  1.135 1.035 1.365 1.295 ;
        RECT  1.150 0.460 1.310 0.750 ;
        RECT  0.385 0.590 1.150 0.750 ;
        RECT  0.975 1.035 1.135 2.230 ;
        RECT  0.285 0.590 0.385 1.290 ;
        RECT  0.285 2.025 0.385 2.285 ;
        RECT  0.225 0.590 0.285 2.285 ;
        RECT  0.125 1.030 0.225 2.285 ;
    END
END SDFFSRHQX2

MACRO SDFFSRHQX1
    CLASS CORE ;
    FOREIGN SDFFSRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.975 1.330 6.315 2.150 ;
        END
        ANTENNAGATEAREA     0.1365 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.820 1.290 5.040 1.845 ;
        RECT  4.725 1.290 4.820 1.580 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 2.100 4.235 2.540 ;
        RECT  3.135 2.380 4.075 2.540 ;
        RECT  2.975 1.290 3.135 2.540 ;
        RECT  2.885 1.290 2.975 1.580 ;
        RECT  2.355 2.380 2.975 2.540 ;
        RECT  2.195 2.165 2.355 2.540 ;
        END
        ANTENNAGATEAREA     0.1261 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.880 1.635 12.140 1.895 ;
        RECT  11.810 1.685 11.880 1.895 ;
        RECT  10.475 1.685 11.810 1.845 ;
        RECT  10.245 1.300 10.475 1.990 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.975 1.290 15.055 2.175 ;
        RECT  14.715 1.035 14.975 2.555 ;
        END
        ANTENNADIFFAREA     0.3944 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.315 1.290 3.555 1.860 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.180 0.435 1.845 ;
        END
        ANTENNAGATEAREA     0.1456 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.425 -0.250 15.180 0.250 ;
        RECT  14.165 -0.250 14.425 0.405 ;
        RECT  12.825 -0.250 14.165 0.250 ;
        RECT  12.565 -0.250 12.825 0.405 ;
        RECT  10.305 -0.250 12.565 0.250 ;
        RECT  10.045 -0.250 10.305 0.405 ;
        RECT  8.700 -0.250 10.045 0.250 ;
        RECT  8.440 -0.250 8.700 0.405 ;
        RECT  5.045 -0.250 8.440 0.250 ;
        RECT  4.785 -0.250 5.045 0.405 ;
        RECT  3.205 -0.250 4.785 0.250 ;
        RECT  2.945 -0.250 3.205 0.405 ;
        RECT  0.895 -0.250 2.945 0.250 ;
        RECT  0.635 -0.250 0.895 0.405 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.425 3.440 15.180 3.940 ;
        RECT  13.825 2.880 14.425 3.940 ;
        RECT  12.435 3.440 13.825 3.940 ;
        RECT  12.175 3.285 12.435 3.940 ;
        RECT  9.155 3.440 12.175 3.940 ;
        RECT  8.895 3.285 9.155 3.940 ;
        RECT  7.755 3.440 8.895 3.940 ;
        RECT  7.495 3.285 7.755 3.940 ;
        RECT  5.635 3.440 7.495 3.940 ;
        RECT  5.375 3.285 5.635 3.940 ;
        RECT  1.235 3.440 5.375 3.940 ;
        RECT  0.635 3.285 1.235 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.205 0.625 14.365 2.695 ;
        RECT  13.515 0.625 14.205 0.785 ;
        RECT  14.105 1.515 14.205 1.775 ;
        RECT  12.945 2.535 14.205 2.695 ;
        RECT  13.895 1.035 13.995 1.295 ;
        RECT  13.895 1.955 13.995 2.215 ;
        RECT  13.735 1.035 13.895 2.215 ;
        RECT  13.535 1.445 13.735 1.705 ;
        RECT  13.255 0.525 13.515 0.785 ;
        RECT  13.215 0.965 13.315 1.225 ;
        RECT  13.215 1.755 13.315 2.015 ;
        RECT  11.630 0.625 13.255 0.785 ;
        RECT  13.055 0.965 13.215 2.355 ;
        RECT  11.305 2.195 13.055 2.355 ;
        RECT  12.685 2.535 12.945 3.155 ;
        RECT  12.735 1.755 12.835 2.015 ;
        RECT  12.575 1.295 12.735 2.015 ;
        RECT  11.645 2.535 12.685 2.695 ;
        RECT  11.190 1.295 12.575 1.455 ;
        RECT  11.485 2.535 11.645 2.810 ;
        RECT  11.470 0.625 11.630 1.065 ;
        RECT  11.370 0.805 11.470 1.065 ;
        RECT  11.145 2.195 11.305 2.760 ;
        RECT  11.030 0.455 11.190 1.455 ;
        RECT  8.555 2.600 11.145 2.760 ;
        RECT  11.085 2.950 11.135 3.210 ;
        RECT  10.875 2.945 11.085 3.210 ;
        RECT  10.840 0.455 11.030 0.745 ;
        RECT  10.705 2.160 10.965 2.420 ;
        RECT  8.465 2.945 10.875 3.105 ;
        RECT  10.690 0.925 10.850 1.205 ;
        RECT  8.260 0.585 10.840 0.745 ;
        RECT  9.335 2.260 10.705 2.420 ;
        RECT  9.435 0.925 10.690 1.085 ;
        RECT  9.335 0.925 9.435 1.185 ;
        RECT  9.175 0.925 9.335 2.420 ;
        RECT  8.735 2.160 9.175 2.420 ;
        RECT  8.835 0.925 8.995 1.980 ;
        RECT  7.915 0.925 8.835 1.085 ;
        RECT  8.555 1.820 8.835 1.980 ;
        RECT  8.305 1.380 8.565 1.640 ;
        RECT  8.395 1.820 8.555 2.760 ;
        RECT  8.205 2.945 8.465 3.250 ;
        RECT  7.575 1.480 8.305 1.640 ;
        RECT  8.100 0.470 8.260 0.745 ;
        RECT  8.055 2.500 8.215 2.760 ;
        RECT  6.655 2.945 8.205 3.105 ;
        RECT  5.385 0.470 8.100 0.630 ;
        RECT  7.445 2.550 8.055 2.760 ;
        RECT  7.755 0.810 7.915 1.085 ;
        RECT  5.795 0.810 7.755 0.970 ;
        RECT  7.445 1.150 7.575 1.640 ;
        RECT  7.285 1.150 7.445 2.760 ;
        RECT  6.835 2.110 7.285 2.370 ;
        RECT  6.655 1.250 6.895 1.510 ;
        RECT  6.495 1.250 6.655 3.260 ;
        RECT  5.975 3.100 6.495 3.260 ;
        RECT  6.155 2.605 6.315 2.920 ;
        RECT  5.385 2.605 6.155 2.765 ;
        RECT  5.815 2.945 5.975 3.260 ;
        RECT  4.915 2.945 5.815 3.105 ;
        RECT  5.635 0.810 5.795 2.190 ;
        RECT  5.565 0.925 5.635 1.185 ;
        RECT  5.225 0.470 5.385 0.745 ;
        RECT  5.225 0.950 5.385 2.765 ;
        RECT  3.270 0.585 5.225 0.745 ;
        RECT  4.090 0.950 5.225 1.110 ;
        RECT  4.755 2.505 5.225 2.765 ;
        RECT  4.885 2.065 5.045 2.325 ;
        RECT  4.755 2.945 4.915 3.220 ;
        RECT  4.575 2.165 4.885 2.325 ;
        RECT  1.675 3.060 4.755 3.220 ;
        RECT  4.415 1.760 4.575 2.880 ;
        RECT  4.235 1.760 4.415 1.920 ;
        RECT  2.015 2.720 4.415 2.880 ;
        RECT  4.075 1.365 4.235 1.920 ;
        RECT  3.735 0.950 3.895 2.200 ;
        RECT  3.495 0.950 3.735 1.110 ;
        RECT  3.485 2.040 3.735 2.200 ;
        RECT  3.110 0.585 3.270 0.930 ;
        RECT  2.775 0.770 3.110 0.930 ;
        RECT  2.695 2.040 2.795 2.200 ;
        RECT  2.695 0.770 2.775 1.110 ;
        RECT  2.535 0.770 2.695 2.200 ;
        RECT  2.515 0.770 2.535 1.110 ;
        RECT  1.620 0.770 2.515 0.930 ;
        RECT  2.015 1.120 2.265 1.280 ;
        RECT  1.280 0.430 2.055 0.590 ;
        RECT  1.855 1.120 2.015 2.880 ;
        RECT  1.515 2.025 1.675 3.220 ;
        RECT  1.460 0.770 1.620 1.845 ;
        RECT  1.115 2.025 1.515 2.185 ;
        RECT  1.295 1.585 1.460 1.845 ;
        RECT  1.120 0.430 1.280 0.810 ;
        RECT  1.115 1.030 1.275 1.290 ;
        RECT  0.775 0.650 1.120 0.810 ;
        RECT  0.955 1.130 1.115 2.185 ;
        RECT  0.615 0.650 0.775 2.200 ;
        RECT  0.385 0.650 0.615 0.810 ;
        RECT  0.385 2.040 0.615 2.200 ;
        RECT  0.125 0.550 0.385 0.810 ;
        RECT  0.225 2.040 0.385 2.770 ;
        RECT  0.125 2.510 0.225 2.770 ;
    END
END SDFFSRHQX1

MACRO SDFFSHQX8
    CLASS CORE ;
    FOREIGN SDFFSHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.780 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.880 1.700 11.375 2.085 ;
        END
        ANTENNAGATEAREA     0.3510 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 1.565 6.775 2.215 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.270 2.225 1.530 ;
        RECT  1.675 1.270 2.175 1.580 ;
        END
        ANTENNAGATEAREA     0.2821 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.820 0.695 19.080 2.895 ;
        RECT  18.060 1.700 18.820 2.400 ;
        RECT  17.800 0.865 18.060 2.895 ;
        END
        ANTENNADIFFAREA     1.5900 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.605 1.505 3.765 1.765 ;
        RECT  3.095 1.505 3.605 1.665 ;
        RECT  2.910 1.290 3.095 1.665 ;
        RECT  2.885 1.290 2.910 1.580 ;
        END
        ANTENNAGATEAREA     0.3016 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.625 0.370 2.190 ;
        END
        ANTENNAGATEAREA     0.4576 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.590 -0.250 19.780 0.250 ;
        RECT  19.330 -0.250 19.590 1.195 ;
        RECT  18.570 -0.250 19.330 0.250 ;
        RECT  18.310 -0.250 18.570 1.095 ;
        RECT  17.660 -0.250 18.310 0.250 ;
        RECT  17.400 -0.250 17.660 0.405 ;
        RECT  15.520 -0.250 17.400 0.250 ;
        RECT  15.880 1.000 16.140 1.260 ;
        RECT  15.520 1.000 15.880 1.160 ;
        RECT  15.360 -0.250 15.520 1.160 ;
        RECT  13.200 -0.250 15.360 0.250 ;
        RECT  12.940 -0.250 13.200 0.575 ;
        RECT  12.115 -0.250 12.940 0.250 ;
        RECT  11.855 -0.250 12.115 0.575 ;
        RECT  11.545 -0.250 11.855 0.250 ;
        RECT  11.285 -0.250 11.545 0.575 ;
        RECT  10.445 -0.250 11.285 0.250 ;
        RECT  10.185 -0.250 10.445 0.625 ;
        RECT  7.250 -0.250 10.185 0.250 ;
        RECT  6.990 -0.250 7.250 0.405 ;
        RECT  5.575 -0.250 6.990 0.250 ;
        RECT  5.315 -0.250 5.575 0.405 ;
        RECT  2.965 -0.250 5.315 0.250 ;
        RECT  2.365 -0.250 2.965 0.405 ;
        RECT  0.385 -0.250 2.365 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.590 3.440 19.780 3.940 ;
        RECT  19.330 1.960 19.590 3.940 ;
        RECT  18.570 3.440 19.330 3.940 ;
        RECT  18.310 2.615 18.570 3.940 ;
        RECT  17.340 3.440 18.310 3.940 ;
        RECT  17.080 3.285 17.340 3.940 ;
        RECT  15.110 3.440 17.080 3.940 ;
        RECT  14.850 3.285 15.110 3.940 ;
        RECT  12.505 3.440 14.850 3.940 ;
        RECT  12.245 2.955 12.505 3.940 ;
        RECT  10.895 3.440 12.245 3.940 ;
        RECT  10.635 3.285 10.895 3.940 ;
        RECT  9.825 3.440 10.635 3.940 ;
        RECT  9.565 3.285 9.825 3.940 ;
        RECT  7.840 3.440 9.565 3.940 ;
        RECT  7.580 3.285 7.840 3.940 ;
        RECT  6.760 3.440 7.580 3.940 ;
        RECT  6.500 3.285 6.760 3.940 ;
        RECT  4.800 3.440 6.500 3.940 ;
        RECT  4.540 3.110 4.800 3.940 ;
        RECT  3.860 3.440 4.540 3.940 ;
        RECT  3.600 3.115 3.860 3.940 ;
        RECT  1.755 3.440 3.600 3.940 ;
        RECT  1.495 3.285 1.755 3.940 ;
        RECT  0.385 3.440 1.495 3.940 ;
        RECT  0.125 2.615 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.460 1.565 17.620 3.105 ;
        RECT  17.395 1.565 17.460 1.725 ;
        RECT  16.720 2.945 17.460 3.105 ;
        RECT  17.235 0.590 17.395 1.725 ;
        RECT  17.120 1.905 17.280 2.750 ;
        RECT  17.220 0.590 17.235 0.750 ;
        RECT  17.060 0.470 17.220 0.750 ;
        RECT  17.000 1.905 17.120 2.065 ;
        RECT  16.300 2.590 17.120 2.750 ;
        RECT  16.140 0.470 17.060 0.630 ;
        RECT  16.880 0.930 17.000 2.065 ;
        RECT  16.660 2.245 16.940 2.405 ;
        RECT  16.840 0.810 16.880 2.065 ;
        RECT  16.620 0.810 16.840 1.090 ;
        RECT  16.510 2.945 16.720 3.260 ;
        RECT  16.500 1.270 16.660 2.405 ;
        RECT  16.010 3.100 16.510 3.260 ;
        RECT  15.525 1.765 16.500 1.925 ;
        RECT  16.140 2.590 16.300 2.865 ;
        RECT  15.880 0.470 16.140 0.750 ;
        RECT  14.845 2.705 16.140 2.865 ;
        RECT  15.700 2.265 15.960 2.525 ;
        RECT  15.185 2.265 15.700 2.425 ;
        RECT  15.365 1.765 15.525 2.045 ;
        RECT  15.125 1.705 15.185 2.425 ;
        RECT  15.025 0.470 15.125 2.425 ;
        RECT  14.965 0.470 15.025 1.865 ;
        RECT  13.540 0.470 14.965 0.630 ;
        RECT  14.780 2.045 14.845 2.865 ;
        RECT  14.685 0.810 14.780 2.865 ;
        RECT  14.620 0.810 14.685 2.205 ;
        RECT  13.880 0.810 14.620 0.970 ;
        RECT  14.045 2.045 14.620 2.205 ;
        RECT  14.345 2.385 14.505 2.985 ;
        RECT  13.565 2.825 14.345 2.985 ;
        RECT  14.220 1.155 14.320 1.315 ;
        RECT  14.060 1.155 14.220 1.725 ;
        RECT  13.565 1.565 14.060 1.725 ;
        RECT  13.785 2.045 14.045 2.645 ;
        RECT  13.720 0.810 13.880 1.315 ;
        RECT  13.425 1.155 13.720 1.315 ;
        RECT  13.405 1.565 13.565 2.985 ;
        RECT  13.425 0.470 13.540 0.915 ;
        RECT  13.380 0.470 13.425 0.945 ;
        RECT  12.875 2.165 13.405 2.425 ;
        RECT  13.165 0.755 13.380 0.945 ;
        RECT  13.065 2.610 13.225 3.215 ;
        RECT  11.005 0.755 13.165 0.915 ;
        RECT  11.790 2.610 13.065 2.775 ;
        RECT  12.715 1.115 12.875 2.425 ;
        RECT  12.395 1.115 12.715 1.275 ;
        RECT  11.995 2.265 12.715 2.425 ;
        RECT  12.225 1.590 12.485 1.850 ;
        RECT  11.715 1.590 12.225 1.750 ;
        RECT  11.735 2.165 11.995 2.425 ;
        RECT  11.630 2.610 11.790 3.105 ;
        RECT  10.665 2.265 11.735 2.425 ;
        RECT  11.555 1.145 11.715 1.750 ;
        RECT  11.625 2.615 11.630 3.105 ;
        RECT  8.400 2.945 11.625 3.105 ;
        RECT  10.215 1.145 11.555 1.305 ;
        RECT  10.215 2.605 11.445 2.765 ;
        RECT  10.955 0.475 11.005 0.915 ;
        RECT  10.745 0.475 10.955 0.965 ;
        RECT  9.355 0.805 10.745 0.965 ;
        RECT  10.505 1.680 10.665 2.425 ;
        RECT  10.405 1.680 10.505 1.940 ;
        RECT  10.055 1.145 10.215 2.765 ;
        RECT  8.870 1.265 10.055 1.425 ;
        RECT  9.925 2.505 10.055 2.765 ;
        RECT  8.845 2.605 9.925 2.765 ;
        RECT  9.715 1.740 9.875 2.250 ;
        RECT  8.400 1.740 9.715 1.900 ;
        RECT  9.190 0.805 9.355 1.085 ;
        RECT  7.645 0.925 9.190 1.085 ;
        RECT  8.585 2.505 8.845 2.765 ;
        RECT  8.240 1.425 8.400 3.105 ;
        RECT  6.255 0.585 8.360 0.745 ;
        RECT  8.100 1.425 8.240 1.685 ;
        RECT  3.010 2.760 8.240 2.920 ;
        RECT  7.865 1.985 8.025 2.245 ;
        RECT  7.645 1.985 7.865 2.145 ;
        RECT  7.485 0.925 7.645 2.145 ;
        RECT  7.200 0.925 7.485 1.085 ;
        RECT  7.200 2.320 7.300 2.580 ;
        RECT  7.040 0.925 7.200 2.580 ;
        RECT  6.435 0.925 7.040 1.085 ;
        RECT  3.350 2.420 7.040 2.580 ;
        RECT  6.255 1.240 6.310 2.180 ;
        RECT  6.150 0.585 6.255 2.180 ;
        RECT  6.095 0.585 6.150 1.400 ;
        RECT  5.620 2.020 6.150 2.180 ;
        RECT  4.785 1.240 6.095 1.400 ;
        RECT  5.810 1.580 5.970 1.840 ;
        RECT  5.755 0.435 5.915 0.745 ;
        RECT  4.545 1.680 5.810 1.840 ;
        RECT  4.785 0.585 5.755 0.745 ;
        RECT  4.105 2.080 5.370 2.240 ;
        RECT  4.625 0.470 4.785 0.745 ;
        RECT  4.625 1.035 4.785 1.400 ;
        RECT  3.325 0.470 4.625 0.630 ;
        RECT  4.445 1.580 4.545 1.840 ;
        RECT  4.285 0.815 4.445 1.840 ;
        RECT  3.665 0.815 4.285 0.975 ;
        RECT  3.945 1.155 4.105 2.240 ;
        RECT  3.845 1.155 3.945 1.315 ;
        RECT  3.570 2.080 3.945 2.240 ;
        RECT  3.505 0.815 3.665 1.085 ;
        RECT  1.745 0.925 3.505 1.085 ;
        RECT  3.190 1.845 3.350 2.580 ;
        RECT  3.165 0.470 3.325 0.745 ;
        RECT  2.665 3.100 3.285 3.260 ;
        RECT  2.705 1.845 3.190 2.005 ;
        RECT  2.085 0.585 3.165 0.745 ;
        RECT  2.850 2.185 3.010 2.920 ;
        RECT  2.205 2.185 2.850 2.345 ;
        RECT  2.505 1.585 2.705 2.005 ;
        RECT  2.505 2.595 2.665 3.260 ;
        RECT  2.445 1.585 2.505 1.845 ;
        RECT  1.865 2.595 2.505 2.755 ;
        RECT  2.165 2.935 2.325 3.195 ;
        RECT  2.045 1.760 2.205 2.345 ;
        RECT  0.895 2.935 2.165 3.095 ;
        RECT  1.925 0.470 2.085 0.745 ;
        RECT  1.405 1.760 2.045 1.920 ;
        RECT  0.725 0.470 1.925 0.630 ;
        RECT  1.705 2.105 1.865 2.755 ;
        RECT  1.585 0.810 1.745 1.085 ;
        RECT  1.065 2.105 1.705 2.265 ;
        RECT  1.065 0.810 1.585 0.970 ;
        RECT  1.245 1.150 1.405 1.920 ;
        RECT  1.035 2.445 1.295 2.705 ;
        RECT  0.905 0.810 1.065 2.265 ;
        RECT  0.725 2.445 1.035 2.605 ;
        RECT  0.635 2.935 0.895 3.215 ;
        RECT  0.565 0.470 0.725 2.605 ;
        RECT  0.125 1.035 0.565 1.295 ;
    END
END SDFFSHQX8

MACRO SDFFSHQX4
    CLASS CORE ;
    FOREIGN SDFFSHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.860 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.880 1.700 11.375 2.085 ;
        END
        ANTENNAGATEAREA     0.3510 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 1.565 6.775 2.215 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.675 1.270 2.175 1.580 ;
        END
        ANTENNAGATEAREA     0.2821 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.965 0.680 18.275 2.895 ;
        END
        ANTENNADIFFAREA     0.8132 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.605 1.505 3.765 1.765 ;
        RECT  3.095 1.505 3.605 1.665 ;
        RECT  2.910 1.290 3.095 1.665 ;
        RECT  2.885 1.290 2.910 1.580 ;
        END
        ANTENNAGATEAREA     0.3016 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.625 0.370 2.190 ;
        END
        ANTENNAGATEAREA     0.4576 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.735 -0.250 18.860 0.250 ;
        RECT  18.475 -0.250 18.735 1.095 ;
        RECT  17.660 -0.250 18.475 0.250 ;
        RECT  17.400 -0.250 17.660 0.405 ;
        RECT  15.520 -0.250 17.400 0.250 ;
        RECT  15.880 1.000 16.140 1.260 ;
        RECT  15.520 1.000 15.880 1.160 ;
        RECT  15.360 -0.250 15.520 1.160 ;
        RECT  13.200 -0.250 15.360 0.250 ;
        RECT  12.940 -0.250 13.200 0.575 ;
        RECT  12.115 -0.250 12.940 0.250 ;
        RECT  11.855 -0.250 12.115 0.575 ;
        RECT  11.545 -0.250 11.855 0.250 ;
        RECT  11.285 -0.250 11.545 0.575 ;
        RECT  10.445 -0.250 11.285 0.250 ;
        RECT  10.185 -0.250 10.445 0.625 ;
        RECT  7.250 -0.250 10.185 0.250 ;
        RECT  6.990 -0.250 7.250 0.405 ;
        RECT  5.575 -0.250 6.990 0.250 ;
        RECT  5.315 -0.250 5.575 0.405 ;
        RECT  2.930 -0.250 5.315 0.250 ;
        RECT  2.330 -0.250 2.930 0.405 ;
        RECT  0.385 -0.250 2.330 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.735 3.440 18.860 3.940 ;
        RECT  18.475 2.275 18.735 3.940 ;
        RECT  17.560 3.440 18.475 3.940 ;
        RECT  17.300 3.285 17.560 3.940 ;
        RECT  15.110 3.440 17.300 3.940 ;
        RECT  14.850 3.285 15.110 3.940 ;
        RECT  12.505 3.440 14.850 3.940 ;
        RECT  12.245 2.955 12.505 3.940 ;
        RECT  10.895 3.440 12.245 3.940 ;
        RECT  10.635 3.285 10.895 3.940 ;
        RECT  9.825 3.440 10.635 3.940 ;
        RECT  9.565 3.285 9.825 3.940 ;
        RECT  7.840 3.440 9.565 3.940 ;
        RECT  7.580 3.285 7.840 3.940 ;
        RECT  6.760 3.440 7.580 3.940 ;
        RECT  6.500 3.285 6.760 3.940 ;
        RECT  4.800 3.440 6.500 3.940 ;
        RECT  4.540 3.110 4.800 3.940 ;
        RECT  3.860 3.440 4.540 3.940 ;
        RECT  3.600 3.115 3.860 3.940 ;
        RECT  1.795 3.440 3.600 3.940 ;
        RECT  1.535 3.285 1.795 3.940 ;
        RECT  0.385 3.440 1.535 3.940 ;
        RECT  0.125 2.615 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.585 0.590 17.745 3.105 ;
        RECT  17.220 0.590 17.585 0.750 ;
        RECT  16.740 2.945 17.585 3.105 ;
        RECT  17.245 1.740 17.405 2.750 ;
        RECT  17.000 1.740 17.245 1.900 ;
        RECT  16.300 2.590 17.245 2.750 ;
        RECT  17.060 0.470 17.220 0.750 ;
        RECT  16.660 2.245 17.065 2.405 ;
        RECT  15.880 0.470 17.060 0.630 ;
        RECT  16.880 0.930 17.000 1.900 ;
        RECT  16.840 0.810 16.880 1.900 ;
        RECT  16.720 0.810 16.840 1.090 ;
        RECT  16.580 2.945 16.740 3.260 ;
        RECT  16.620 0.810 16.720 0.970 ;
        RECT  16.500 1.270 16.660 2.405 ;
        RECT  16.135 3.100 16.580 3.260 ;
        RECT  15.525 1.765 16.500 1.925 ;
        RECT  16.140 2.590 16.300 2.865 ;
        RECT  14.845 2.705 16.140 2.865 ;
        RECT  15.700 2.265 15.960 2.525 ;
        RECT  15.185 2.265 15.700 2.425 ;
        RECT  15.365 1.765 15.525 2.045 ;
        RECT  15.120 1.705 15.185 2.425 ;
        RECT  15.025 0.470 15.120 2.425 ;
        RECT  14.960 0.470 15.025 1.865 ;
        RECT  13.540 0.470 14.960 0.630 ;
        RECT  14.780 2.045 14.845 2.865 ;
        RECT  14.685 0.810 14.780 2.865 ;
        RECT  14.620 0.810 14.685 2.205 ;
        RECT  13.880 0.810 14.620 0.970 ;
        RECT  14.045 2.045 14.620 2.205 ;
        RECT  14.345 2.385 14.505 2.985 ;
        RECT  13.565 2.825 14.345 2.985 ;
        RECT  14.220 1.155 14.320 1.315 ;
        RECT  14.060 1.155 14.220 1.725 ;
        RECT  13.565 1.565 14.060 1.725 ;
        RECT  13.785 2.045 14.045 2.645 ;
        RECT  13.720 0.810 13.880 1.315 ;
        RECT  13.425 1.155 13.720 1.315 ;
        RECT  13.405 1.565 13.565 2.985 ;
        RECT  13.425 0.470 13.540 0.915 ;
        RECT  13.380 0.470 13.425 0.945 ;
        RECT  12.875 2.165 13.405 2.425 ;
        RECT  13.165 0.755 13.380 0.945 ;
        RECT  13.065 2.615 13.225 3.215 ;
        RECT  11.005 0.755 13.165 0.915 ;
        RECT  11.795 2.615 13.065 2.775 ;
        RECT  12.715 1.115 12.875 2.425 ;
        RECT  12.395 1.115 12.715 1.275 ;
        RECT  11.995 2.265 12.715 2.425 ;
        RECT  12.225 1.590 12.485 1.850 ;
        RECT  11.715 1.590 12.225 1.750 ;
        RECT  11.735 2.165 11.995 2.425 ;
        RECT  11.635 2.615 11.795 3.105 ;
        RECT  10.665 2.265 11.735 2.425 ;
        RECT  11.555 1.145 11.715 1.750 ;
        RECT  8.405 2.945 11.635 3.105 ;
        RECT  10.215 1.145 11.555 1.305 ;
        RECT  10.215 2.605 11.445 2.765 ;
        RECT  10.955 0.475 11.005 0.915 ;
        RECT  10.745 0.475 10.955 0.965 ;
        RECT  9.355 0.805 10.745 0.965 ;
        RECT  10.505 1.680 10.665 2.425 ;
        RECT  10.405 1.680 10.505 1.940 ;
        RECT  10.055 1.145 10.215 2.765 ;
        RECT  8.870 1.265 10.055 1.425 ;
        RECT  9.925 2.505 10.055 2.765 ;
        RECT  8.845 2.605 9.925 2.765 ;
        RECT  9.715 1.740 9.875 2.250 ;
        RECT  8.405 1.740 9.715 1.900 ;
        RECT  9.190 0.805 9.355 1.085 ;
        RECT  7.645 0.925 9.190 1.085 ;
        RECT  8.585 2.505 8.845 2.765 ;
        RECT  8.245 1.420 8.405 3.105 ;
        RECT  6.255 0.585 8.360 0.745 ;
        RECT  8.150 1.420 8.245 1.685 ;
        RECT  3.010 2.760 8.245 2.920 ;
        RECT  8.100 1.425 8.150 1.685 ;
        RECT  7.865 1.985 8.025 2.245 ;
        RECT  7.645 1.985 7.865 2.145 ;
        RECT  7.485 0.925 7.645 2.145 ;
        RECT  7.175 0.925 7.485 1.085 ;
        RECT  7.175 2.320 7.300 2.580 ;
        RECT  7.015 0.925 7.175 2.580 ;
        RECT  6.435 0.925 7.015 1.085 ;
        RECT  3.350 2.420 7.015 2.580 ;
        RECT  6.255 1.240 6.310 2.240 ;
        RECT  6.150 0.585 6.255 2.240 ;
        RECT  6.095 0.585 6.150 1.400 ;
        RECT  5.620 2.080 6.150 2.240 ;
        RECT  4.785 1.240 6.095 1.400 ;
        RECT  5.810 1.580 5.970 1.840 ;
        RECT  5.755 0.435 5.915 0.745 ;
        RECT  4.545 1.680 5.810 1.840 ;
        RECT  4.785 0.585 5.755 0.745 ;
        RECT  4.105 2.080 5.370 2.240 ;
        RECT  4.625 0.470 4.785 0.745 ;
        RECT  4.625 1.035 4.785 1.400 ;
        RECT  3.285 0.470 4.625 0.630 ;
        RECT  4.445 1.580 4.545 1.840 ;
        RECT  4.285 0.815 4.445 1.840 ;
        RECT  3.625 0.815 4.285 0.975 ;
        RECT  3.945 1.155 4.105 2.240 ;
        RECT  3.810 1.155 3.945 1.315 ;
        RECT  3.570 2.080 3.945 2.240 ;
        RECT  3.465 0.815 3.625 1.085 ;
        RECT  1.745 0.925 3.465 1.085 ;
        RECT  3.190 1.845 3.350 2.580 ;
        RECT  3.125 0.470 3.285 0.745 ;
        RECT  2.665 3.100 3.285 3.260 ;
        RECT  2.665 1.845 3.190 2.005 ;
        RECT  2.085 0.585 3.125 0.745 ;
        RECT  2.850 2.185 3.010 2.920 ;
        RECT  2.180 2.185 2.850 2.345 ;
        RECT  2.505 1.585 2.665 2.005 ;
        RECT  2.505 2.595 2.665 3.260 ;
        RECT  2.405 1.585 2.505 1.845 ;
        RECT  1.830 2.595 2.505 2.755 ;
        RECT  2.165 2.935 2.325 3.195 ;
        RECT  2.020 1.760 2.180 2.345 ;
        RECT  0.895 2.935 2.165 3.095 ;
        RECT  1.925 0.470 2.085 0.745 ;
        RECT  1.405 1.760 2.020 1.920 ;
        RECT  0.725 0.470 1.925 0.630 ;
        RECT  1.670 2.105 1.830 2.755 ;
        RECT  1.585 0.810 1.745 1.085 ;
        RECT  1.065 2.105 1.670 2.265 ;
        RECT  1.065 0.810 1.585 0.970 ;
        RECT  1.245 1.150 1.405 1.920 ;
        RECT  1.035 2.445 1.295 2.705 ;
        RECT  0.905 0.810 1.065 2.265 ;
        RECT  0.725 2.445 1.035 2.605 ;
        RECT  0.635 2.935 0.895 3.215 ;
        RECT  0.565 0.470 0.725 2.605 ;
        RECT  0.125 1.035 0.565 1.295 ;
    END
END SDFFSHQX4

MACRO SDFFSHQX2
    CLASS CORE ;
    FOREIGN SDFFSHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.800 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.285 1.630 8.340 2.085 ;
        RECT  8.025 1.575 8.285 2.085 ;
        RECT  7.945 1.630 8.025 2.085 ;
        END
        ANTENNAGATEAREA     0.2054 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.585 1.625 5.010 1.990 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.880 1.290 2.225 1.665 ;
        END
        ANTENNAGATEAREA     0.1755 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.235 0.695 13.390 1.295 ;
        RECT  13.075 0.695 13.235 2.600 ;
        RECT  13.005 1.515 13.075 2.600 ;
        RECT  12.975 2.000 13.005 2.600 ;
        END
        ANTENNADIFFAREA     0.5668 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.845 2.710 2.195 ;
        RECT  2.425 1.700 2.635 2.195 ;
        RECT  2.340 1.845 2.425 2.195 ;
        END
        ANTENNAGATEAREA     0.1703 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.475 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2626 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.850 -0.250 13.800 0.250 ;
        RECT  12.590 -0.250 12.850 1.050 ;
        RECT  10.375 -0.250 12.590 0.250 ;
        RECT  10.115 -0.250 10.375 0.405 ;
        RECT  8.585 -0.250 10.115 0.250 ;
        RECT  8.325 -0.250 8.585 0.405 ;
        RECT  7.960 -0.250 8.325 0.250 ;
        RECT  7.800 -0.250 7.960 0.655 ;
        RECT  5.490 -0.250 7.800 0.250 ;
        RECT  5.230 -0.250 5.490 0.405 ;
        RECT  4.550 -0.250 5.230 0.250 ;
        RECT  4.290 -0.250 4.550 0.405 ;
        RECT  2.595 -0.250 4.290 0.250 ;
        RECT  2.335 -0.250 2.595 0.405 ;
        RECT  0.335 -0.250 2.335 0.250 ;
        RECT  0.175 -0.250 0.335 0.640 ;
        RECT  0.000 -0.250 0.175 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.635 3.440 13.800 3.940 ;
        RECT  13.035 3.060 13.635 3.940 ;
        RECT  10.395 3.440 13.035 3.940 ;
        RECT  10.135 3.065 10.395 3.940 ;
        RECT  8.845 3.440 10.135 3.940 ;
        RECT  8.585 3.115 8.845 3.940 ;
        RECT  7.245 3.440 8.585 3.940 ;
        RECT  6.985 3.285 7.245 3.940 ;
        RECT  5.625 3.440 6.985 3.940 ;
        RECT  5.365 2.905 5.625 3.940 ;
        RECT  4.715 3.440 5.365 3.940 ;
        RECT  4.455 3.285 4.715 3.940 ;
        RECT  2.390 3.440 4.455 3.940 ;
        RECT  2.230 3.060 2.390 3.940 ;
        RECT  0.860 3.440 2.230 3.940 ;
        RECT  0.600 2.890 0.860 3.940 ;
        RECT  0.000 3.440 0.600 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.635 1.230 12.795 3.165 ;
        RECT  12.410 1.230 12.635 1.390 ;
        RECT  12.235 3.005 12.635 3.165 ;
        RECT  12.295 1.575 12.455 2.825 ;
        RECT  12.250 0.430 12.410 1.390 ;
        RECT  12.195 1.575 12.295 1.835 ;
        RECT  11.725 2.665 12.295 2.825 ;
        RECT  11.625 0.430 12.250 0.590 ;
        RECT  11.560 3.005 12.235 3.235 ;
        RECT  12.065 1.575 12.195 1.735 ;
        RECT  11.950 2.000 12.110 2.270 ;
        RECT  11.905 0.770 12.065 1.735 ;
        RECT  11.430 2.000 11.950 2.170 ;
        RECT  11.805 0.770 11.905 0.930 ;
        RECT  11.465 2.630 11.725 2.825 ;
        RECT  11.465 0.430 11.625 0.695 ;
        RECT  10.955 0.525 11.465 0.695 ;
        RECT  10.695 2.665 11.465 2.825 ;
        RECT  11.270 1.035 11.430 2.170 ;
        RECT  11.170 1.035 11.270 1.485 ;
        RECT  10.745 1.325 11.170 1.485 ;
        RECT  10.875 1.665 11.035 2.465 ;
        RECT  10.695 0.525 10.955 0.795 ;
        RECT  10.235 1.665 10.875 1.825 ;
        RECT  10.485 1.225 10.745 1.485 ;
        RECT  10.535 2.045 10.695 2.825 ;
        RECT  9.895 2.045 10.535 2.205 ;
        RECT  10.195 2.385 10.355 2.645 ;
        RECT  10.075 0.585 10.235 1.825 ;
        RECT  9.385 2.435 10.195 2.595 ;
        RECT  9.895 0.585 10.075 0.745 ;
        RECT  9.635 0.430 9.895 0.745 ;
        RECT  9.795 1.995 9.895 2.255 ;
        RECT  9.635 1.065 9.795 2.255 ;
        RECT  9.385 2.775 9.645 3.095 ;
        RECT  8.300 0.585 9.635 0.745 ;
        RECT  9.375 0.965 9.635 1.225 ;
        RECT  9.125 2.310 9.385 2.595 ;
        RECT  8.135 2.775 9.385 2.935 ;
        RECT  8.965 0.960 9.125 2.595 ;
        RECT  8.865 0.960 8.965 1.220 ;
        RECT  8.205 2.435 8.965 2.595 ;
        RECT  8.680 1.400 8.780 2.000 ;
        RECT  8.520 1.175 8.680 2.000 ;
        RECT  7.845 1.175 8.520 1.335 ;
        RECT  8.140 0.585 8.300 0.995 ;
        RECT  8.045 2.265 8.205 2.595 ;
        RECT  7.590 0.835 8.140 0.995 ;
        RECT  7.975 2.775 8.135 3.105 ;
        RECT  7.030 2.265 8.045 2.425 ;
        RECT  6.705 2.945 7.975 3.105 ;
        RECT  7.685 1.175 7.845 1.445 ;
        RECT  6.690 2.605 7.795 2.765 ;
        RECT  6.690 1.285 7.685 1.445 ;
        RECT  7.505 0.475 7.590 0.995 ;
        RECT  7.340 0.475 7.505 1.105 ;
        RECT  6.350 0.945 7.340 1.105 ;
        RECT  6.900 0.475 7.160 0.745 ;
        RECT  6.870 1.710 7.030 2.425 ;
        RECT  6.005 0.585 6.900 0.745 ;
        RECT  6.445 2.945 6.705 3.205 ;
        RECT  6.530 1.285 6.690 2.765 ;
        RECT  6.235 2.325 6.530 2.765 ;
        RECT  6.055 2.945 6.445 3.105 ;
        RECT  6.190 0.945 6.350 1.425 ;
        RECT  6.055 1.615 6.200 1.875 ;
        RECT  5.715 1.265 6.190 1.425 ;
        RECT  5.895 1.615 6.055 3.105 ;
        RECT  5.845 0.585 6.005 1.085 ;
        RECT  5.090 2.565 5.895 2.725 ;
        RECT  4.405 0.925 5.845 1.085 ;
        RECT  5.555 1.265 5.715 2.385 ;
        RECT  4.800 1.265 5.555 1.425 ;
        RECT  4.745 2.225 5.555 2.385 ;
        RECT  4.930 2.565 5.090 3.105 ;
        RECT  4.840 0.435 5.000 0.745 ;
        RECT  2.730 2.945 4.930 3.105 ;
        RECT  2.135 0.585 4.840 0.745 ;
        RECT  4.585 2.225 4.745 2.765 ;
        RECT  3.075 2.605 4.585 2.765 ;
        RECT  4.245 0.925 4.405 2.425 ;
        RECT  3.760 1.135 4.245 1.295 ;
        RECT  3.715 2.265 4.245 2.425 ;
        RECT  3.905 1.795 4.065 2.055 ;
        RECT  3.830 1.795 3.905 1.955 ;
        RECT  3.670 1.655 3.830 1.955 ;
        RECT  3.600 0.930 3.760 1.295 ;
        RECT  3.390 1.655 3.670 1.815 ;
        RECT  3.255 1.995 3.415 2.425 ;
        RECT  3.230 0.925 3.390 1.815 ;
        RECT  3.050 1.995 3.255 2.155 ;
        RECT  1.965 0.925 3.230 1.085 ;
        RECT  2.915 2.375 3.075 2.765 ;
        RECT  2.890 1.265 3.050 2.155 ;
        RECT  2.160 2.375 2.915 2.535 ;
        RECT  2.765 1.265 2.890 1.425 ;
        RECT  2.570 2.715 2.730 3.105 ;
        RECT  1.790 2.715 2.570 2.875 ;
        RECT  2.000 1.845 2.160 2.535 ;
        RECT  1.975 0.480 2.135 0.745 ;
        RECT  1.695 1.845 2.000 2.005 ;
        RECT  0.675 0.480 1.975 0.640 ;
        RECT  1.795 0.925 1.965 1.105 ;
        RECT  1.230 3.055 1.870 3.215 ;
        RECT  1.635 0.825 1.795 1.105 ;
        RECT  1.630 2.185 1.790 2.875 ;
        RECT  1.535 1.655 1.695 2.005 ;
        RECT  1.015 0.825 1.635 0.985 ;
        RECT  1.355 2.185 1.630 2.345 ;
        RECT  1.355 1.165 1.455 1.325 ;
        RECT  1.195 1.165 1.355 2.345 ;
        RECT  1.070 2.525 1.230 3.215 ;
        RECT  1.015 2.525 1.070 2.685 ;
        RECT  0.855 0.825 1.015 2.685 ;
        RECT  0.515 0.480 0.675 2.345 ;
        RECT  0.200 1.035 0.515 1.295 ;
        RECT  0.460 2.185 0.515 2.345 ;
        RECT  0.200 2.185 0.460 2.445 ;
    END
END SDFFSHQX2

MACRO SDFFSHQX1
    CLASS CORE ;
    FOREIGN SDFFSHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.420 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.405 1.700 8.615 1.990 ;
        RECT  7.825 1.705 8.405 1.865 ;
        END
        ANTENNAGATEAREA     0.1352 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.775 1.630 4.935 2.070 ;
        RECT  4.615 1.625 4.775 2.070 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.265 2.175 1.580 ;
        RECT  1.630 1.265 1.965 1.550 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.395 1.700 11.655 2.215 ;
        RECT  11.375 1.700 11.395 1.990 ;
        RECT  11.325 1.105 11.375 1.990 ;
        RECT  11.165 0.985 11.325 1.990 ;
        RECT  11.105 0.985 11.165 1.245 ;
        END
        ANTENNADIFFAREA     0.3460 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.700 2.635 2.105 ;
        RECT  2.270 1.780 2.425 2.105 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.475 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1560 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.815 -0.250 12.420 0.250 ;
        RECT  11.655 -0.250 11.815 0.810 ;
        RECT  10.075 -0.250 11.655 0.250 ;
        RECT  9.815 -0.250 10.075 0.405 ;
        RECT  8.405 -0.250 9.815 0.250 ;
        RECT  8.145 -0.250 8.405 0.405 ;
        RECT  7.770 -0.250 8.145 0.250 ;
        RECT  7.510 -0.250 7.770 0.655 ;
        RECT  5.380 -0.250 7.510 0.250 ;
        RECT  5.120 -0.250 5.380 0.405 ;
        RECT  4.475 -0.250 5.120 0.250 ;
        RECT  4.215 -0.250 4.475 0.405 ;
        RECT  2.345 -0.250 4.215 0.250 ;
        RECT  2.085 -0.250 2.345 0.405 ;
        RECT  0.815 -0.250 2.085 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.995 3.440 12.420 3.940 ;
        RECT  11.735 3.075 11.995 3.940 ;
        RECT  7.830 3.440 11.735 3.940 ;
        RECT  7.570 3.115 7.830 3.940 ;
        RECT  7.125 3.440 7.570 3.940 ;
        RECT  6.865 3.285 7.125 3.940 ;
        RECT  5.315 3.440 6.865 3.940 ;
        RECT  5.055 3.285 5.315 3.940 ;
        RECT  4.405 3.440 5.055 3.940 ;
        RECT  4.145 3.285 4.405 3.940 ;
        RECT  2.085 3.440 4.145 3.940 ;
        RECT  1.925 3.015 2.085 3.940 ;
        RECT  0.815 3.440 1.925 3.940 ;
        RECT  0.555 2.890 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.185 1.035 12.295 1.295 ;
        RECT  12.025 0.430 12.185 1.295 ;
        RECT  11.995 2.480 12.065 2.740 ;
        RECT  11.995 1.135 12.025 1.295 ;
        RECT  11.835 1.135 11.995 2.740 ;
        RECT  11.805 2.480 11.835 2.740 ;
        RECT  11.340 2.480 11.805 2.640 ;
        RECT  11.180 2.480 11.340 3.165 ;
        RECT  9.905 3.005 11.180 3.165 ;
        RECT  10.925 1.485 10.985 2.640 ;
        RECT  10.825 0.575 10.925 2.640 ;
        RECT  10.765 0.575 10.825 1.690 ;
        RECT  9.295 2.480 10.825 2.640 ;
        RECT  10.735 0.575 10.765 0.735 ;
        RECT  10.475 0.475 10.735 0.735 ;
        RECT  10.585 1.905 10.625 2.165 ;
        RECT  10.425 0.985 10.585 2.165 ;
        RECT  10.400 1.725 10.425 2.165 ;
        RECT  10.045 1.725 10.400 1.985 ;
        RECT  9.475 0.580 9.635 2.295 ;
        RECT  9.345 3.005 9.605 3.220 ;
        RECT  9.060 0.580 9.475 0.740 ;
        RECT  8.175 3.060 9.345 3.220 ;
        RECT  9.135 0.920 9.295 2.770 ;
        RECT  9.105 0.920 9.135 1.180 ;
        RECT  8.975 2.510 9.135 2.770 ;
        RECT  8.955 0.450 9.060 0.740 ;
        RECT  8.795 0.450 8.955 0.745 ;
        RECT  8.925 1.360 8.955 2.330 ;
        RECT  8.795 0.925 8.925 2.330 ;
        RECT  8.110 0.585 8.795 0.745 ;
        RECT  8.765 0.925 8.795 1.520 ;
        RECT  8.725 2.170 8.795 2.330 ;
        RECT  8.545 0.925 8.765 1.085 ;
        RECT  8.465 2.170 8.725 2.875 ;
        RECT  8.375 1.360 8.565 1.520 ;
        RECT  8.045 2.170 8.465 2.330 ;
        RECT  8.215 1.285 8.375 1.520 ;
        RECT  6.545 1.285 8.215 1.445 ;
        RECT  8.010 2.770 8.175 3.220 ;
        RECT  7.950 0.585 8.110 0.995 ;
        RECT  7.885 2.045 8.045 2.330 ;
        RECT  6.800 2.770 8.010 2.930 ;
        RECT  7.295 0.835 7.950 0.995 ;
        RECT  7.605 2.045 7.885 2.205 ;
        RECT  6.545 2.385 7.705 2.545 ;
        RECT  7.445 1.625 7.605 2.205 ;
        RECT  7.345 1.625 7.445 1.785 ;
        RECT  7.230 0.475 7.295 0.995 ;
        RECT  7.035 0.475 7.230 1.105 ;
        RECT  7.030 0.525 7.035 1.105 ;
        RECT  5.480 0.945 7.030 1.105 ;
        RECT  6.555 0.475 6.815 0.745 ;
        RECT  6.640 2.770 6.800 3.105 ;
        RECT  6.630 2.945 6.640 3.105 ;
        RECT  6.370 2.945 6.630 3.115 ;
        RECT  5.140 0.585 6.555 0.745 ;
        RECT  6.385 1.285 6.545 2.545 ;
        RECT  6.175 2.275 6.385 2.545 ;
        RECT  5.990 2.945 6.370 3.105 ;
        RECT  5.845 1.585 5.990 3.105 ;
        RECT  5.830 1.535 5.845 3.105 ;
        RECT  5.685 1.535 5.830 1.795 ;
        RECT  2.425 2.945 5.830 3.105 ;
        RECT  5.490 2.015 5.650 2.665 ;
        RECT  4.915 2.505 5.490 2.665 ;
        RECT  5.320 0.945 5.480 1.425 ;
        RECT  4.435 1.265 5.320 1.425 ;
        RECT  4.980 0.585 5.140 1.085 ;
        RECT  4.095 0.925 4.980 1.085 ;
        RECT  4.435 2.505 4.915 2.765 ;
        RECT  4.640 0.485 4.800 0.745 ;
        RECT  0.675 0.585 4.640 0.745 ;
        RECT  4.275 1.265 4.435 2.765 ;
        RECT  2.765 2.605 4.275 2.765 ;
        RECT  3.935 0.925 4.095 2.425 ;
        RECT  3.685 1.135 3.935 1.295 ;
        RECT  3.405 2.265 3.935 2.425 ;
        RECT  3.595 1.520 3.755 2.055 ;
        RECT  3.525 0.925 3.685 1.295 ;
        RECT  3.315 1.520 3.595 1.680 ;
        RECT  3.155 0.925 3.315 1.680 ;
        RECT  1.015 0.925 3.155 1.085 ;
        RECT  2.975 1.910 3.105 2.425 ;
        RECT  2.945 1.265 2.975 2.425 ;
        RECT  2.815 1.265 2.945 2.070 ;
        RECT  2.690 1.265 2.815 1.425 ;
        RECT  2.605 2.335 2.765 2.765 ;
        RECT  2.085 2.335 2.605 2.495 ;
        RECT  2.265 2.675 2.425 3.105 ;
        RECT  1.745 2.675 2.265 2.835 ;
        RECT  1.925 1.845 2.085 2.495 ;
        RECT  1.695 1.845 1.925 2.005 ;
        RECT  1.585 2.185 1.745 2.835 ;
        RECT  1.535 1.745 1.695 2.005 ;
        RECT  1.355 2.185 1.585 2.345 ;
        RECT  1.395 3.055 1.565 3.215 ;
        RECT  1.235 2.525 1.395 3.215 ;
        RECT  1.195 1.265 1.355 2.345 ;
        RECT  1.015 2.525 1.235 2.685 ;
        RECT  0.855 0.925 1.015 2.685 ;
        RECT  0.515 0.585 0.675 2.345 ;
        RECT  0.125 1.035 0.515 1.295 ;
        RECT  0.385 2.185 0.515 2.345 ;
        RECT  0.125 2.185 0.385 2.445 ;
    END
END SDFFSHQX1

MACRO SDFFRHQX8
    CLASS CORE ;
    FOREIGN SDFFRHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.275 5.460 1.775 ;
        END
        ANTENNAGATEAREA     0.1534 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.225 1.835 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.040 1.885 13.200 2.145 ;
        RECT  10.915 1.985 13.040 2.145 ;
        RECT  10.915 1.275 10.950 1.535 ;
        RECT  10.705 1.275 10.915 2.145 ;
        RECT  9.700 1.275 10.705 1.435 ;
        RECT  10.580 1.855 10.705 2.145 ;
        RECT  10.425 1.855 10.580 2.115 ;
        RECT  9.440 1.275 9.700 1.535 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.760 1.515 16.895 1.765 ;
        RECT  16.500 0.600 16.760 3.055 ;
        RECT  15.740 1.300 16.500 2.400 ;
        RECT  15.480 0.600 15.740 3.055 ;
        RECT  15.305 1.220 15.480 3.055 ;
        END
        ANTENNADIFFAREA     1.6264 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.655 2.705 1.915 ;
        RECT  2.475 1.290 2.635 1.915 ;
        RECT  2.425 1.290 2.475 1.580 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.545 0.625 1.990 ;
        END
        ANTENNAGATEAREA     0.3744 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.270 -0.250 17.480 0.250 ;
        RECT  17.010 -0.250 17.270 1.095 ;
        RECT  16.250 -0.250 17.010 0.250 ;
        RECT  15.990 -0.250 16.250 1.120 ;
        RECT  15.200 -0.250 15.990 0.250 ;
        RECT  14.940 -0.250 15.200 0.840 ;
        RECT  13.990 -0.250 14.940 0.250 ;
        RECT  13.730 -0.250 13.990 0.405 ;
        RECT  11.320 -0.250 13.730 0.250 ;
        RECT  11.060 -0.250 11.320 0.405 ;
        RECT  9.455 -0.250 11.060 0.250 ;
        RECT  9.195 -0.250 9.455 0.405 ;
        RECT  8.350 -0.250 9.195 0.250 ;
        RECT  8.090 -0.250 8.350 0.405 ;
        RECT  6.590 -0.250 8.090 0.250 ;
        RECT  6.430 -0.250 6.590 0.935 ;
        RECT  4.845 -0.250 6.430 0.250 ;
        RECT  4.585 -0.250 4.845 0.405 ;
        RECT  1.955 -0.250 4.585 0.250 ;
        RECT  1.695 -0.250 1.955 0.405 ;
        RECT  0.815 -0.250 1.695 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.270 3.440 17.480 3.940 ;
        RECT  17.010 2.275 17.270 3.940 ;
        RECT  16.250 3.440 17.010 3.940 ;
        RECT  15.990 2.615 16.250 3.940 ;
        RECT  15.040 3.440 15.990 3.940 ;
        RECT  14.780 2.955 15.040 3.940 ;
        RECT  13.630 3.440 14.780 3.940 ;
        RECT  13.370 3.065 13.630 3.940 ;
        RECT  10.260 3.440 13.370 3.940 ;
        RECT  10.000 3.285 10.260 3.940 ;
        RECT  9.160 3.440 10.000 3.940 ;
        RECT  8.900 3.285 9.160 3.940 ;
        RECT  7.905 3.440 8.900 3.940 ;
        RECT  7.645 2.945 7.905 3.940 ;
        RECT  6.170 3.440 7.645 3.940 ;
        RECT  5.910 3.285 6.170 3.940 ;
        RECT  5.220 3.440 5.910 3.940 ;
        RECT  4.960 3.285 5.220 3.940 ;
        RECT  2.825 3.440 4.960 3.940 ;
        RECT  2.565 3.115 2.825 3.940 ;
        RECT  0.725 3.440 2.565 3.940 ;
        RECT  0.125 2.845 0.725 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.015 1.545 15.115 1.805 ;
        RECT  14.855 1.545 15.015 2.775 ;
        RECT  14.435 2.615 14.855 2.775 ;
        RECT  14.560 1.955 14.660 2.215 ;
        RECT  14.400 1.035 14.560 2.215 ;
        RECT  14.175 2.615 14.435 2.880 ;
        RECT  14.060 0.585 14.220 2.435 ;
        RECT  13.880 2.665 14.175 2.825 ;
        RECT  12.060 0.585 14.060 0.745 ;
        RECT  13.720 0.925 13.880 2.825 ;
        RECT  11.630 0.925 13.720 1.085 ;
        RECT  12.415 2.665 13.720 2.825 ;
        RECT  13.380 1.365 13.540 2.485 ;
        RECT  12.260 1.365 13.380 1.525 ;
        RECT  11.905 2.325 13.380 2.485 ;
        RECT  12.925 3.005 13.185 3.220 ;
        RECT  10.630 3.060 12.925 3.220 ;
        RECT  12.185 2.665 12.415 2.880 ;
        RECT  12.000 1.265 12.260 1.525 ;
        RECT  11.135 2.720 12.185 2.880 ;
        RECT  11.800 0.440 12.060 0.745 ;
        RECT  11.290 1.365 12.000 1.525 ;
        RECT  11.740 2.325 11.905 2.540 ;
        RECT  8.910 0.585 11.800 0.745 ;
        RECT  10.885 2.380 11.740 2.540 ;
        RECT  11.470 0.925 11.630 1.185 ;
        RECT  11.130 0.925 11.290 1.525 ;
        RECT  10.090 0.925 11.130 1.085 ;
        RECT  10.625 2.380 10.885 2.715 ;
        RECT  10.470 2.945 10.630 3.220 ;
        RECT  9.710 2.380 10.625 2.540 ;
        RECT  8.460 2.945 10.470 3.105 ;
        RECT  9.945 1.635 10.205 1.880 ;
        RECT  9.230 1.720 9.945 1.880 ;
        RECT  9.450 2.165 9.710 2.765 ;
        RECT  8.890 2.380 9.450 2.540 ;
        RECT  9.070 1.085 9.230 1.880 ;
        RECT  8.480 1.085 9.070 1.245 ;
        RECT  8.650 0.510 8.910 0.905 ;
        RECT  8.730 1.430 8.890 2.540 ;
        RECT  6.940 0.745 8.650 0.905 ;
        RECT  8.320 1.085 8.480 2.275 ;
        RECT  8.300 2.560 8.460 3.105 ;
        RECT  7.230 1.085 8.320 1.245 ;
        RECT  8.265 2.115 8.320 2.275 ;
        RECT  8.200 2.560 8.300 2.820 ;
        RECT  8.005 2.115 8.265 2.380 ;
        RECT  7.375 2.560 8.200 2.720 ;
        RECT  8.040 1.460 8.140 1.620 ;
        RECT  7.880 1.460 8.040 1.870 ;
        RECT  7.035 2.115 8.005 2.275 ;
        RECT  6.840 1.710 7.880 1.870 ;
        RECT  7.215 2.560 7.375 3.055 ;
        RECT  6.595 2.895 7.215 3.055 ;
        RECT  6.775 2.115 7.035 2.715 ;
        RECT  6.780 0.745 6.940 1.275 ;
        RECT  6.595 1.455 6.840 1.870 ;
        RECT  6.200 1.115 6.780 1.275 ;
        RECT  6.580 1.455 6.595 3.055 ;
        RECT  6.435 1.710 6.580 3.055 ;
        RECT  3.225 2.895 6.435 3.055 ;
        RECT  6.060 0.455 6.220 0.775 ;
        RECT  6.040 0.955 6.200 2.255 ;
        RECT  5.530 0.615 6.060 0.775 ;
        RECT  5.750 0.955 6.040 1.115 ;
        RECT  5.770 2.095 6.040 2.255 ;
        RECT  5.510 2.095 5.770 2.715 ;
        RECT  5.370 0.615 5.530 1.085 ;
        RECT  3.565 2.555 5.510 2.715 ;
        RECT  4.970 0.925 5.370 1.085 ;
        RECT  5.025 0.480 5.185 0.745 ;
        RECT  4.100 0.585 5.025 0.745 ;
        RECT  4.810 0.925 4.970 2.185 ;
        RECT  3.755 0.925 4.810 1.085 ;
        RECT  4.510 2.025 4.810 2.185 ;
        RECT  4.470 1.455 4.630 1.845 ;
        RECT  4.350 2.025 4.510 2.370 ;
        RECT  3.415 1.455 4.470 1.615 ;
        RECT  4.250 2.110 4.350 2.370 ;
        RECT  3.940 0.480 4.100 0.745 ;
        RECT  3.740 2.095 4.000 2.375 ;
        RECT  2.295 0.480 3.940 0.640 ;
        RECT  3.595 0.825 3.755 1.085 ;
        RECT  3.075 2.095 3.740 2.255 ;
        RECT  3.405 2.435 3.565 2.715 ;
        RECT  3.255 0.820 3.415 1.615 ;
        RECT  1.675 2.435 3.405 2.595 ;
        RECT  2.635 0.820 3.255 0.980 ;
        RECT  3.065 2.775 3.225 3.055 ;
        RECT  2.915 1.160 3.075 2.255 ;
        RECT  1.675 2.775 3.065 2.935 ;
        RECT  2.815 1.160 2.915 1.320 ;
        RECT  2.755 2.095 2.915 2.255 ;
        RECT  2.475 0.820 2.635 1.085 ;
        RECT  1.785 0.925 2.475 1.085 ;
        RECT  2.135 0.480 2.295 0.745 ;
        RECT  0.965 0.585 2.135 0.745 ;
        RECT  1.785 2.020 2.075 2.180 ;
        RECT  1.625 0.925 1.785 2.180 ;
        RECT  1.445 2.775 1.675 3.035 ;
        RECT  1.415 1.025 1.445 3.035 ;
        RECT  1.405 1.025 1.415 2.935 ;
        RECT  1.285 0.930 1.405 2.935 ;
        RECT  1.145 0.930 1.285 1.190 ;
        RECT  0.805 0.585 0.965 2.345 ;
        RECT  0.125 0.905 0.805 1.165 ;
        RECT  0.385 2.185 0.805 2.345 ;
        RECT  0.125 2.185 0.385 2.445 ;
    END
END SDFFRHQX8

MACRO SDFFRHQX4
    CLASS CORE ;
    FOREIGN SDFFRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.560 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.275 5.460 1.775 ;
        END
        ANTENNAGATEAREA     0.1534 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.225 1.835 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.040 1.885 13.200 2.145 ;
        RECT  10.890 1.985 13.040 2.145 ;
        RECT  10.915 1.275 10.950 1.535 ;
        RECT  10.890 1.275 10.915 1.700 ;
        RECT  10.790 1.275 10.890 2.145 ;
        RECT  10.705 1.290 10.790 2.145 ;
        RECT  9.700 1.295 10.705 1.455 ;
        RECT  10.475 1.855 10.705 2.145 ;
        RECT  9.440 1.275 9.700 1.535 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.695 2.115 15.740 3.055 ;
        RECT  15.480 0.645 15.695 3.055 ;
        RECT  15.435 0.645 15.480 2.810 ;
        RECT  15.305 1.105 15.435 2.810 ;
        END
        ANTENNADIFFAREA     0.8132 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.655 2.705 1.915 ;
        RECT  2.475 1.290 2.635 1.915 ;
        RECT  2.425 1.290 2.475 1.580 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.545 0.625 1.990 ;
        END
        ANTENNAGATEAREA     0.3744 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.205 -0.250 16.560 0.250 ;
        RECT  15.945 -0.250 16.205 1.120 ;
        RECT  15.110 -0.250 15.945 0.250 ;
        RECT  14.850 -0.250 15.110 0.840 ;
        RECT  13.990 -0.250 14.850 0.250 ;
        RECT  13.730 -0.250 13.990 0.405 ;
        RECT  11.320 -0.250 13.730 0.250 ;
        RECT  11.060 -0.250 11.320 0.405 ;
        RECT  9.455 -0.250 11.060 0.250 ;
        RECT  9.195 -0.250 9.455 0.405 ;
        RECT  8.350 -0.250 9.195 0.250 ;
        RECT  8.090 -0.250 8.350 0.405 ;
        RECT  6.590 -0.250 8.090 0.250 ;
        RECT  6.430 -0.250 6.590 0.935 ;
        RECT  4.845 -0.250 6.430 0.250 ;
        RECT  4.585 -0.250 4.845 0.405 ;
        RECT  1.955 -0.250 4.585 0.250 ;
        RECT  1.695 -0.250 1.955 0.405 ;
        RECT  0.815 -0.250 1.695 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.250 3.440 16.560 3.940 ;
        RECT  15.990 2.170 16.250 3.940 ;
        RECT  15.040 3.440 15.990 3.940 ;
        RECT  14.780 2.955 15.040 3.940 ;
        RECT  13.630 3.440 14.780 3.940 ;
        RECT  13.370 3.065 13.630 3.940 ;
        RECT  10.260 3.440 13.370 3.940 ;
        RECT  10.000 3.285 10.260 3.940 ;
        RECT  9.160 3.440 10.000 3.940 ;
        RECT  8.900 3.285 9.160 3.940 ;
        RECT  7.905 3.440 8.900 3.940 ;
        RECT  7.645 2.945 7.905 3.940 ;
        RECT  6.170 3.440 7.645 3.940 ;
        RECT  5.910 3.285 6.170 3.940 ;
        RECT  5.220 3.440 5.910 3.940 ;
        RECT  4.960 3.285 5.220 3.940 ;
        RECT  2.825 3.440 4.960 3.940 ;
        RECT  2.565 3.115 2.825 3.940 ;
        RECT  0.725 3.440 2.565 3.940 ;
        RECT  0.125 2.825 0.725 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.085 1.545 15.115 1.805 ;
        RECT  14.925 1.545 15.085 2.775 ;
        RECT  14.855 1.545 14.925 1.805 ;
        RECT  14.435 2.615 14.925 2.775 ;
        RECT  14.560 1.955 14.675 2.215 ;
        RECT  14.400 1.035 14.560 2.215 ;
        RECT  14.175 2.615 14.435 2.880 ;
        RECT  14.060 0.585 14.220 2.435 ;
        RECT  13.880 2.665 14.175 2.825 ;
        RECT  12.060 0.585 14.060 0.745 ;
        RECT  13.720 0.925 13.880 2.825 ;
        RECT  12.800 0.925 13.720 1.085 ;
        RECT  12.415 2.665 13.720 2.825 ;
        RECT  13.380 1.365 13.540 2.485 ;
        RECT  12.260 1.365 13.380 1.525 ;
        RECT  11.905 2.325 13.380 2.485 ;
        RECT  12.925 3.005 13.185 3.220 ;
        RECT  10.630 3.060 12.925 3.220 ;
        RECT  12.540 0.925 12.800 1.185 ;
        RECT  11.630 0.925 12.540 1.085 ;
        RECT  12.145 2.665 12.415 2.880 ;
        RECT  12.000 1.265 12.260 1.525 ;
        RECT  11.135 2.720 12.145 2.880 ;
        RECT  11.800 0.440 12.060 0.745 ;
        RECT  11.290 1.365 12.000 1.525 ;
        RECT  11.625 2.325 11.905 2.540 ;
        RECT  8.910 0.585 11.800 0.745 ;
        RECT  11.470 0.925 11.630 1.185 ;
        RECT  10.885 2.380 11.625 2.540 ;
        RECT  11.130 0.925 11.290 1.525 ;
        RECT  10.090 0.925 11.130 1.085 ;
        RECT  10.625 2.380 10.885 2.715 ;
        RECT  10.470 2.945 10.630 3.220 ;
        RECT  9.710 2.380 10.625 2.540 ;
        RECT  8.460 2.945 10.470 3.105 ;
        RECT  9.945 1.635 10.205 1.885 ;
        RECT  9.230 1.725 9.945 1.885 ;
        RECT  9.450 2.070 9.710 2.670 ;
        RECT  8.890 2.070 9.450 2.230 ;
        RECT  9.070 1.085 9.230 1.885 ;
        RECT  8.480 1.085 9.070 1.245 ;
        RECT  8.650 0.510 8.910 0.840 ;
        RECT  8.730 1.430 8.890 2.230 ;
        RECT  6.940 0.680 8.650 0.840 ;
        RECT  8.320 1.085 8.480 2.275 ;
        RECT  8.300 2.560 8.460 3.105 ;
        RECT  7.490 1.085 8.320 1.245 ;
        RECT  8.265 2.115 8.320 2.275 ;
        RECT  8.200 2.560 8.300 2.820 ;
        RECT  8.005 2.115 8.265 2.380 ;
        RECT  7.375 2.560 8.200 2.720 ;
        RECT  8.040 1.425 8.140 1.685 ;
        RECT  7.880 1.425 8.040 1.870 ;
        RECT  7.035 2.115 8.005 2.275 ;
        RECT  6.840 1.710 7.880 1.870 ;
        RECT  7.230 1.035 7.490 1.295 ;
        RECT  7.215 2.560 7.375 3.055 ;
        RECT  6.595 2.895 7.215 3.055 ;
        RECT  6.775 2.115 7.035 2.715 ;
        RECT  6.780 0.680 6.940 1.275 ;
        RECT  6.595 1.455 6.840 1.870 ;
        RECT  6.250 1.115 6.780 1.275 ;
        RECT  6.580 1.455 6.595 3.055 ;
        RECT  6.435 1.710 6.580 3.055 ;
        RECT  3.165 2.895 6.435 3.055 ;
        RECT  6.150 1.115 6.250 1.665 ;
        RECT  6.060 0.455 6.220 0.775 ;
        RECT  5.990 0.955 6.150 2.255 ;
        RECT  5.530 0.615 6.060 0.775 ;
        RECT  5.750 0.955 5.990 1.115 ;
        RECT  5.770 2.095 5.990 2.255 ;
        RECT  5.510 2.095 5.770 2.715 ;
        RECT  5.370 0.615 5.530 1.085 ;
        RECT  3.505 2.555 5.510 2.715 ;
        RECT  4.970 0.925 5.370 1.085 ;
        RECT  5.025 0.480 5.185 0.745 ;
        RECT  4.100 0.585 5.025 0.745 ;
        RECT  4.810 0.925 4.970 2.225 ;
        RECT  3.755 0.925 4.810 1.085 ;
        RECT  4.510 2.065 4.810 2.225 ;
        RECT  4.470 1.405 4.630 1.845 ;
        RECT  4.250 2.065 4.510 2.325 ;
        RECT  3.700 1.405 4.470 1.565 ;
        RECT  3.940 0.480 4.100 0.745 ;
        RECT  3.740 2.095 4.000 2.375 ;
        RECT  2.295 0.480 3.940 0.640 ;
        RECT  3.595 0.825 3.755 1.085 ;
        RECT  3.075 2.095 3.740 2.255 ;
        RECT  3.440 1.405 3.700 1.665 ;
        RECT  3.345 2.435 3.505 2.715 ;
        RECT  3.415 1.405 3.440 1.565 ;
        RECT  3.255 0.820 3.415 1.565 ;
        RECT  1.675 2.435 3.345 2.595 ;
        RECT  2.635 0.820 3.255 0.980 ;
        RECT  3.005 2.775 3.165 3.055 ;
        RECT  2.915 1.160 3.075 2.255 ;
        RECT  1.675 2.775 3.005 2.935 ;
        RECT  2.815 1.160 2.915 1.320 ;
        RECT  2.755 2.095 2.915 2.255 ;
        RECT  2.475 0.820 2.635 1.085 ;
        RECT  1.785 0.925 2.475 1.085 ;
        RECT  2.135 0.480 2.295 0.745 ;
        RECT  0.965 0.585 2.135 0.745 ;
        RECT  1.785 2.020 2.075 2.180 ;
        RECT  1.625 0.925 1.785 2.180 ;
        RECT  1.445 2.775 1.675 3.035 ;
        RECT  1.415 1.035 1.445 3.035 ;
        RECT  1.405 1.035 1.415 2.935 ;
        RECT  1.285 0.965 1.405 2.935 ;
        RECT  1.145 0.965 1.285 1.225 ;
        RECT  0.805 0.585 0.965 2.330 ;
        RECT  0.125 0.905 0.805 1.165 ;
        RECT  0.385 2.170 0.805 2.330 ;
        RECT  0.125 2.170 0.385 2.430 ;
    END
END SDFFRHQX4

MACRO SDFFRHQX2
    CLASS CORE ;
    FOREIGN SDFFRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.420 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.295 4.475 1.990 ;
        RECT  4.230 1.295 4.265 1.565 ;
        END
        ANTENNAGATEAREA     0.0832 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.175 1.580 ;
        RECT  1.540 1.290 1.965 1.530 ;
        END
        ANTENNAGATEAREA     0.1833 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.330 1.605 9.450 1.765 ;
        RECT  9.170 1.605 9.330 1.900 ;
        RECT  9.075 1.700 9.170 1.900 ;
        RECT  8.570 1.740 9.075 1.900 ;
        RECT  8.470 1.740 8.570 2.065 ;
        RECT  8.410 1.740 8.470 2.275 ;
        RECT  8.310 1.805 8.410 2.275 ;
        RECT  7.695 2.115 8.310 2.275 ;
        RECT  7.645 1.700 7.695 2.275 ;
        RECT  7.535 1.510 7.645 2.275 ;
        RECT  7.485 1.510 7.535 1.990 ;
        RECT  7.330 1.510 7.485 1.670 ;
        END
        ANTENNAGATEAREA     0.2366 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.270 1.515 12.295 2.995 ;
        RECT  12.170 1.515 12.270 3.055 ;
        RECT  12.010 1.035 12.170 3.055 ;
        RECT  11.995 1.035 12.010 1.195 ;
        RECT  11.735 0.595 11.995 1.195 ;
        END
        ANTENNADIFFAREA     0.7276 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 1.635 2.635 2.090 ;
        END
        ANTENNAGATEAREA     0.1586 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.475 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2444 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.420 -0.250 12.420 0.250 ;
        RECT  11.160 -0.250 11.420 0.840 ;
        RECT  9.890 -0.250 11.160 0.250 ;
        RECT  9.630 -0.250 9.890 0.405 ;
        RECT  7.235 -0.250 9.630 0.250 ;
        RECT  6.975 -0.250 7.235 0.405 ;
        RECT  5.355 -0.250 6.975 0.250 ;
        RECT  5.095 -0.250 5.355 0.405 ;
        RECT  4.475 -0.250 5.095 0.250 ;
        RECT  4.215 -0.250 4.475 0.405 ;
        RECT  2.495 -0.250 4.215 0.250 ;
        RECT  2.235 -0.250 2.495 0.405 ;
        RECT  0.335 -0.250 2.235 0.250 ;
        RECT  0.175 -0.250 0.335 0.630 ;
        RECT  0.000 -0.250 0.175 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.720 3.440 12.420 3.940 ;
        RECT  11.460 2.955 11.720 3.940 ;
        RECT  10.265 3.440 11.460 3.940 ;
        RECT  10.005 3.065 10.265 3.940 ;
        RECT  8.265 3.440 10.005 3.940 ;
        RECT  8.005 3.285 8.265 3.940 ;
        RECT  7.325 3.440 8.005 3.940 ;
        RECT  7.065 3.285 7.325 3.940 ;
        RECT  5.580 3.440 7.065 3.940 ;
        RECT  5.320 3.285 5.580 3.940 ;
        RECT  4.640 3.440 5.320 3.940 ;
        RECT  4.380 3.285 4.640 3.940 ;
        RECT  2.350 3.440 4.380 3.940 ;
        RECT  2.190 2.950 2.350 3.940 ;
        RECT  0.815 3.440 2.190 3.940 ;
        RECT  0.555 2.895 0.815 3.940 ;
        RECT  0.215 2.895 0.555 3.155 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.655 1.545 11.755 1.805 ;
        RECT  11.495 1.545 11.655 2.760 ;
        RECT  11.005 2.600 11.495 2.760 ;
        RECT  11.215 1.955 11.300 2.215 ;
        RECT  11.200 1.530 11.215 2.215 ;
        RECT  11.040 1.525 11.200 2.215 ;
        RECT  10.865 1.525 11.040 1.690 ;
        RECT  10.745 2.600 11.005 2.965 ;
        RECT  10.705 1.035 10.865 1.690 ;
        RECT  10.545 2.105 10.805 2.365 ;
        RECT  10.185 2.600 10.745 2.760 ;
        RECT  10.525 2.105 10.545 2.265 ;
        RECT  10.365 0.585 10.525 2.265 ;
        RECT  9.235 0.585 10.365 0.745 ;
        RECT  10.025 0.925 10.185 2.760 ;
        RECT  8.720 0.925 10.025 1.085 ;
        RECT  9.095 2.600 10.025 2.760 ;
        RECT  9.685 1.265 9.845 2.415 ;
        RECT  8.380 1.265 9.685 1.425 ;
        RECT  8.860 2.255 9.685 2.415 ;
        RECT  8.805 3.005 9.525 3.165 ;
        RECT  9.075 0.470 9.235 0.745 ;
        RECT  8.580 0.470 9.075 0.630 ;
        RECT  8.700 2.255 8.860 2.715 ;
        RECT  8.645 2.945 8.805 3.165 ;
        RECT  8.560 0.825 8.720 1.085 ;
        RECT  8.585 2.455 8.700 2.715 ;
        RECT  5.800 2.945 8.645 3.105 ;
        RECT  7.865 2.455 8.585 2.615 ;
        RECT  8.320 0.440 8.580 0.630 ;
        RECT  8.220 0.815 8.380 1.425 ;
        RECT  7.575 0.470 8.320 0.630 ;
        RECT  7.980 0.815 8.220 0.975 ;
        RECT  7.880 1.155 8.040 1.935 ;
        RECT  6.380 1.155 7.880 1.315 ;
        RECT  7.605 2.455 7.865 2.715 ;
        RECT  7.110 2.455 7.605 2.615 ;
        RECT  7.415 0.470 7.575 0.970 ;
        RECT  6.735 0.810 7.415 0.970 ;
        RECT  6.950 1.800 7.110 2.615 ;
        RECT  6.850 1.800 6.950 2.060 ;
        RECT  6.475 0.430 6.735 0.970 ;
        RECT  6.035 0.805 6.475 0.970 ;
        RECT  6.380 2.440 6.430 2.700 ;
        RECT  6.220 1.155 6.380 2.700 ;
        RECT  5.695 0.465 6.255 0.625 ;
        RECT  6.170 2.440 6.220 2.700 ;
        RECT  5.875 0.805 6.035 1.425 ;
        RECT  5.155 1.265 5.875 1.425 ;
        RECT  5.640 1.605 5.800 3.105 ;
        RECT  5.535 0.465 5.695 1.085 ;
        RECT  5.540 1.605 5.640 1.765 ;
        RECT  2.690 2.945 5.640 3.105 ;
        RECT  4.815 0.925 5.535 1.085 ;
        RECT  5.180 1.750 5.270 2.055 ;
        RECT  5.155 1.750 5.180 2.765 ;
        RECT  4.995 1.265 5.155 2.765 ;
        RECT  3.030 2.605 4.995 2.765 ;
        RECT  4.655 0.505 4.915 0.745 ;
        RECT  4.655 0.925 4.815 2.395 ;
        RECT  2.035 0.585 4.655 0.745 ;
        RECT  3.685 0.925 4.655 1.085 ;
        RECT  3.670 2.235 4.655 2.395 ;
        RECT  3.890 1.590 4.050 2.050 ;
        RECT  3.315 1.590 3.890 1.750 ;
        RECT  3.525 0.925 3.685 1.185 ;
        RECT  3.210 1.930 3.370 2.425 ;
        RECT  3.155 0.950 3.315 1.750 ;
        RECT  2.975 1.930 3.210 2.090 ;
        RECT  1.695 0.950 3.155 1.110 ;
        RECT  2.870 2.270 3.030 2.765 ;
        RECT  2.815 1.295 2.975 2.090 ;
        RECT  2.135 2.270 2.870 2.430 ;
        RECT  2.690 1.295 2.815 1.455 ;
        RECT  2.530 2.610 2.690 3.105 ;
        RECT  1.795 2.610 2.530 2.770 ;
        RECT  1.975 1.845 2.135 2.430 ;
        RECT  1.875 0.470 2.035 0.745 ;
        RECT  1.695 1.845 1.975 2.005 ;
        RECT  0.675 0.470 1.875 0.630 ;
        RECT  1.155 3.000 1.825 3.160 ;
        RECT  1.635 2.185 1.795 2.770 ;
        RECT  1.535 0.815 1.695 1.110 ;
        RECT  1.535 1.710 1.695 2.005 ;
        RECT  1.535 2.185 1.635 2.445 ;
        RECT  1.015 0.815 1.535 0.975 ;
        RECT  1.355 2.185 1.535 2.345 ;
        RECT  1.195 1.155 1.355 2.345 ;
        RECT  1.015 2.525 1.155 3.160 ;
        RECT  0.995 0.815 1.015 3.160 ;
        RECT  0.855 0.815 0.995 2.685 ;
        RECT  0.515 0.470 0.675 2.345 ;
        RECT  0.125 1.035 0.515 1.295 ;
        RECT  0.385 2.185 0.515 2.345 ;
        RECT  0.125 2.185 0.385 2.445 ;
    END
END SDFFRHQX2

MACRO SDFFRHQX1
    CLASS CORE ;
    FOREIGN SDFFRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.775 1.630 4.935 2.070 ;
        RECT  4.615 1.625 4.775 2.070 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.650 1.290 2.175 1.580 ;
        END
        ANTENNAGATEAREA     0.1274 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.095 1.660 9.255 1.990 ;
        RECT  9.050 1.700 9.095 1.990 ;
        RECT  8.615 1.830 9.050 1.990 ;
        RECT  8.405 1.700 8.615 1.990 ;
        RECT  8.325 1.830 8.405 1.990 ;
        RECT  8.065 1.830 8.325 2.275 ;
        RECT  7.425 1.830 8.065 1.990 ;
        RECT  7.165 1.730 7.425 1.990 ;
        END
        ANTENNAGATEAREA     0.1430 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.800 1.105 11.835 2.400 ;
        RECT  11.795 0.970 11.800 2.400 ;
        RECT  11.640 0.970 11.795 2.580 ;
        RECT  11.625 0.970 11.640 1.765 ;
        RECT  11.535 1.980 11.640 2.580 ;
        RECT  11.540 0.970 11.625 1.230 ;
        END
        ANTENNADIFFAREA     0.3965 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.365 1.700 2.635 2.155 ;
        END
        ANTENNAGATEAREA     0.0897 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.475 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.255 -0.250 11.960 0.250 ;
        RECT  10.995 -0.250 11.255 0.840 ;
        RECT  9.825 -0.250 10.995 0.250 ;
        RECT  9.565 -0.250 9.825 0.405 ;
        RECT  7.175 -0.250 9.565 0.250 ;
        RECT  6.915 -0.250 7.175 0.405 ;
        RECT  5.565 -0.250 6.915 0.250 ;
        RECT  5.305 -0.250 5.565 0.405 ;
        RECT  4.475 -0.250 5.305 0.250 ;
        RECT  4.215 -0.250 4.475 0.405 ;
        RECT  2.345 -0.250 4.215 0.250 ;
        RECT  2.085 -0.250 2.345 0.405 ;
        RECT  0.815 -0.250 2.085 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.245 3.440 11.960 3.940 ;
        RECT  10.985 3.285 11.245 3.940 ;
        RECT  9.680 3.440 10.985 3.940 ;
        RECT  9.420 3.065 9.680 3.940 ;
        RECT  8.075 3.440 9.420 3.940 ;
        RECT  7.815 3.285 8.075 3.940 ;
        RECT  7.225 3.440 7.815 3.940 ;
        RECT  6.965 3.285 7.225 3.940 ;
        RECT  5.455 3.440 6.965 3.940 ;
        RECT  5.195 3.285 5.455 3.940 ;
        RECT  4.405 3.440 5.195 3.940 ;
        RECT  4.145 3.285 4.405 3.940 ;
        RECT  2.085 3.440 4.145 3.940 ;
        RECT  1.925 3.015 2.085 3.940 ;
        RECT  0.815 3.440 1.925 3.940 ;
        RECT  0.555 2.895 0.815 3.940 ;
        RECT  0.215 2.895 0.555 3.155 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.135 1.485 11.235 1.745 ;
        RECT  10.975 1.485 11.135 2.825 ;
        RECT  10.570 2.665 10.975 2.825 ;
        RECT  10.700 1.035 10.750 1.295 ;
        RECT  10.540 1.035 10.700 2.240 ;
        RECT  10.310 2.665 10.570 3.000 ;
        RECT  10.465 1.035 10.540 1.690 ;
        RECT  10.275 2.220 10.320 2.480 ;
        RECT  9.935 2.665 10.310 2.825 ;
        RECT  10.115 0.585 10.275 2.480 ;
        RECT  9.310 0.585 10.115 0.745 ;
        RECT  9.775 0.925 9.935 2.825 ;
        RECT  8.535 0.925 9.775 1.085 ;
        RECT  9.165 2.665 9.775 2.825 ;
        RECT  9.435 1.265 9.595 2.370 ;
        RECT  8.195 1.265 9.435 1.425 ;
        RECT  8.665 2.210 9.435 2.370 ;
        RECT  9.150 0.470 9.310 0.745 ;
        RECT  8.905 2.550 9.165 2.825 ;
        RECT  8.800 0.470 9.150 0.630 ;
        RECT  8.540 0.445 8.800 0.630 ;
        RECT  8.555 2.945 8.715 3.215 ;
        RECT  8.505 2.210 8.665 2.715 ;
        RECT  5.990 2.945 8.555 3.105 ;
        RECT  7.540 0.470 8.540 0.630 ;
        RECT  8.375 0.810 8.535 1.085 ;
        RECT  8.395 2.455 8.505 2.715 ;
        RECT  7.675 2.455 8.395 2.615 ;
        RECT  8.035 0.910 8.195 1.425 ;
        RECT  7.775 0.810 8.035 1.070 ;
        RECT  7.695 1.285 7.855 1.545 ;
        RECT  6.335 1.285 7.695 1.445 ;
        RECT  7.415 2.455 7.675 2.715 ;
        RECT  7.380 0.470 7.540 1.085 ;
        RECT  6.945 2.455 7.415 2.615 ;
        RECT  6.635 0.925 7.380 1.085 ;
        RECT  6.785 1.625 6.945 2.615 ;
        RECT  6.685 1.625 6.785 1.785 ;
        RECT  6.375 0.650 6.635 1.085 ;
        RECT  5.880 0.925 6.375 1.085 ;
        RECT  6.175 1.285 6.335 2.525 ;
        RECT  6.170 1.285 6.175 1.445 ;
        RECT  5.885 0.485 6.145 0.745 ;
        RECT  5.830 1.705 5.990 3.105 ;
        RECT  5.540 0.585 5.885 0.745 ;
        RECT  5.720 0.925 5.880 1.425 ;
        RECT  5.665 1.705 5.830 1.865 ;
        RECT  2.425 2.945 5.830 3.105 ;
        RECT  4.435 1.265 5.720 1.425 ;
        RECT  5.405 1.605 5.665 1.865 ;
        RECT  5.490 2.085 5.650 2.665 ;
        RECT  5.380 0.585 5.540 1.085 ;
        RECT  4.915 2.505 5.490 2.665 ;
        RECT  4.095 0.925 5.380 1.085 ;
        RECT  4.860 0.485 5.120 0.745 ;
        RECT  4.435 2.505 4.915 2.765 ;
        RECT  0.675 0.585 4.860 0.745 ;
        RECT  4.275 1.265 4.435 2.765 ;
        RECT  2.765 2.605 4.275 2.765 ;
        RECT  3.935 0.925 4.095 2.425 ;
        RECT  3.685 1.135 3.935 1.295 ;
        RECT  3.405 2.265 3.935 2.425 ;
        RECT  3.595 1.655 3.755 2.055 ;
        RECT  3.525 1.035 3.685 1.295 ;
        RECT  3.315 1.655 3.595 1.815 ;
        RECT  3.155 0.925 3.315 1.815 ;
        RECT  1.915 0.925 3.155 1.085 ;
        RECT  2.975 1.995 3.105 2.425 ;
        RECT  2.945 1.265 2.975 2.425 ;
        RECT  2.815 1.265 2.945 2.155 ;
        RECT  2.690 1.265 2.815 1.425 ;
        RECT  2.605 2.335 2.765 2.765 ;
        RECT  2.135 2.335 2.605 2.495 ;
        RECT  2.265 2.675 2.425 3.105 ;
        RECT  1.795 2.675 2.265 2.835 ;
        RECT  1.975 1.860 2.135 2.495 ;
        RECT  1.695 1.860 1.975 2.020 ;
        RECT  1.655 0.925 1.915 1.105 ;
        RECT  1.635 2.200 1.795 2.835 ;
        RECT  1.535 1.760 1.695 2.020 ;
        RECT  1.015 0.925 1.655 1.085 ;
        RECT  1.535 2.200 1.635 2.460 ;
        RECT  1.155 3.055 1.565 3.215 ;
        RECT  1.355 2.200 1.535 2.360 ;
        RECT  1.195 1.265 1.355 2.360 ;
        RECT  1.015 2.540 1.155 3.215 ;
        RECT  0.995 0.925 1.015 3.215 ;
        RECT  0.855 0.925 0.995 2.700 ;
        RECT  0.515 0.585 0.675 2.345 ;
        RECT  0.125 1.035 0.515 1.295 ;
        RECT  0.385 2.185 0.515 2.345 ;
        RECT  0.125 2.185 0.385 2.445 ;
    END
END SDFFRHQX1

MACRO SDFFHQX8
    CLASS CORE ;
    FOREIGN SDFFHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.100 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.085 1.235 5.395 1.990 ;
        END
        ANTENNAGATEAREA     0.1443 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.575 2.225 1.835 ;
        RECT  1.965 1.290 2.175 1.835 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.410 1.515 15.515 1.765 ;
        RECT  15.150 0.595 15.410 3.055 ;
        RECT  14.390 1.700 15.150 2.400 ;
        RECT  14.130 0.595 14.390 3.055 ;
        END
        ANTENNADIFFAREA     1.6264 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.545 2.705 1.915 ;
        RECT  2.545 1.290 2.635 1.915 ;
        RECT  2.450 1.290 2.545 1.705 ;
        RECT  2.425 1.290 2.450 1.580 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.455 0.385 2.015 ;
        END
        ANTENNAGATEAREA     0.3731 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.920 -0.250 16.100 0.250 ;
        RECT  15.660 -0.250 15.920 1.095 ;
        RECT  14.900 -0.250 15.660 0.250 ;
        RECT  14.640 -0.250 14.900 1.095 ;
        RECT  13.880 -0.250 14.640 0.250 ;
        RECT  13.620 -0.250 13.880 0.755 ;
        RECT  12.910 -0.250 13.620 0.250 ;
        RECT  12.650 -0.250 12.910 0.950 ;
        RECT  10.190 -0.250 12.650 0.250 ;
        RECT  9.930 -0.250 10.190 0.405 ;
        RECT  9.250 -0.250 9.930 0.250 ;
        RECT  8.990 -0.250 9.250 0.405 ;
        RECT  8.135 -0.250 8.990 0.250 ;
        RECT  7.875 -0.250 8.135 0.405 ;
        RECT  6.545 -0.250 7.875 0.250 ;
        RECT  6.385 -0.250 6.545 1.070 ;
        RECT  4.985 -0.250 6.385 0.250 ;
        RECT  6.205 0.810 6.385 1.070 ;
        RECT  4.725 -0.250 4.985 0.625 ;
        RECT  1.955 -0.250 4.725 0.250 ;
        RECT  1.695 -0.250 1.955 0.405 ;
        RECT  0.815 -0.250 1.695 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.920 3.440 16.100 3.940 ;
        RECT  15.660 2.275 15.920 3.940 ;
        RECT  14.900 3.440 15.660 3.940 ;
        RECT  14.640 2.615 14.900 3.940 ;
        RECT  13.880 3.440 14.640 3.940 ;
        RECT  13.280 2.955 13.880 3.940 ;
        RECT  10.210 3.440 13.280 3.940 ;
        RECT  9.950 3.285 10.210 3.940 ;
        RECT  9.130 3.440 9.950 3.940 ;
        RECT  8.870 3.285 9.130 3.940 ;
        RECT  7.495 3.440 8.870 3.940 ;
        RECT  7.235 3.285 7.495 3.940 ;
        RECT  6.135 3.440 7.235 3.940 ;
        RECT  5.875 3.285 6.135 3.940 ;
        RECT  5.335 3.440 5.875 3.940 ;
        RECT  5.075 3.285 5.335 3.940 ;
        RECT  3.415 3.440 5.075 3.940 ;
        RECT  2.475 3.115 3.415 3.940 ;
        RECT  0.725 3.440 2.475 3.940 ;
        RECT  0.125 2.805 0.725 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.790 1.510 13.860 1.770 ;
        RECT  13.630 1.510 13.790 2.730 ;
        RECT  13.600 1.510 13.630 1.770 ;
        RECT  12.480 2.570 13.630 2.730 ;
        RECT  13.370 1.035 13.420 1.295 ;
        RECT  13.370 2.040 13.420 2.300 ;
        RECT  13.210 1.035 13.370 2.300 ;
        RECT  13.160 1.035 13.210 1.295 ;
        RECT  12.790 1.500 13.210 1.760 ;
        RECT  13.160 2.040 13.210 2.300 ;
        RECT  12.480 2.065 12.740 2.325 ;
        RECT  12.460 2.065 12.480 2.225 ;
        RECT  12.040 2.505 12.480 2.765 ;
        RECT  12.300 0.470 12.460 2.225 ;
        RECT  12.140 2.960 12.400 3.220 ;
        RECT  10.530 0.470 12.300 0.630 ;
        RECT  10.550 3.060 12.140 3.220 ;
        RECT  11.960 1.200 12.120 1.530 ;
        RECT  11.880 2.165 12.040 2.765 ;
        RECT  11.210 1.200 11.960 1.360 ;
        RECT  11.210 2.165 11.880 2.325 ;
        RECT  10.870 0.810 11.770 0.970 ;
        RECT  11.370 2.505 11.630 2.765 ;
        RECT  10.610 2.605 11.370 2.765 ;
        RECT  11.120 1.150 11.210 2.325 ;
        RECT  11.050 1.150 11.120 2.425 ;
        RECT  10.860 2.165 11.050 2.425 ;
        RECT  10.710 0.810 10.870 1.085 ;
        RECT  10.700 0.925 10.710 1.085 ;
        RECT  10.440 0.925 10.700 1.185 ;
        RECT  10.350 2.485 10.610 2.765 ;
        RECT  10.390 2.945 10.550 3.220 ;
        RECT  10.370 0.470 10.530 0.745 ;
        RECT  9.840 0.925 10.440 1.085 ;
        RECT  8.720 2.945 10.390 3.105 ;
        RECT  7.575 0.585 10.370 0.745 ;
        RECT  9.670 2.605 10.350 2.765 ;
        RECT  9.680 0.925 9.840 2.170 ;
        RECT  9.530 0.925 9.680 1.185 ;
        RECT  9.670 2.010 9.680 2.170 ;
        RECT  9.410 2.010 9.670 2.765 ;
        RECT  9.240 1.515 9.500 1.775 ;
        RECT  8.860 2.010 9.410 2.170 ;
        RECT  9.205 1.515 9.240 1.675 ;
        RECT  9.045 0.955 9.205 1.675 ;
        RECT  8.250 0.955 9.045 1.115 ;
        RECT  8.700 1.535 8.860 2.170 ;
        RECT  8.460 2.845 8.720 3.105 ;
        RECT  8.600 1.535 8.700 1.795 ;
        RECT  6.075 2.945 8.460 3.105 ;
        RECT  8.250 2.405 8.350 2.665 ;
        RECT  8.090 0.955 8.250 2.665 ;
        RECT  7.235 0.955 8.090 1.115 ;
        RECT  6.645 2.505 8.090 2.665 ;
        RECT  7.415 0.470 7.575 0.745 ;
        RECT  7.170 1.905 7.430 2.165 ;
        RECT  6.885 0.470 7.415 0.630 ;
        RECT  7.075 0.905 7.235 1.165 ;
        RECT  6.885 1.905 7.170 2.065 ;
        RECT  6.725 0.470 6.885 2.065 ;
        RECT  5.955 1.250 6.725 1.410 ;
        RECT  6.385 2.490 6.645 2.750 ;
        RECT  6.125 1.590 6.385 1.850 ;
        RECT  5.335 0.470 6.205 0.630 ;
        RECT  6.075 1.690 6.125 1.850 ;
        RECT  5.915 1.690 6.075 3.105 ;
        RECT  5.735 0.865 5.955 1.410 ;
        RECT  4.675 2.945 5.915 3.105 ;
        RECT  5.575 0.865 5.735 2.765 ;
        RECT  5.475 2.215 5.575 2.765 ;
        RECT  1.675 2.435 5.475 2.595 ;
        RECT  5.175 0.470 5.335 0.970 ;
        RECT  4.905 0.810 5.175 0.970 ;
        RECT  4.745 0.810 4.905 2.255 ;
        RECT  4.005 0.810 4.745 0.970 ;
        RECT  4.215 2.095 4.745 2.255 ;
        RECT  4.515 2.775 4.675 3.105 ;
        RECT  4.405 1.585 4.565 1.845 ;
        RECT  1.675 2.775 4.515 2.935 ;
        RECT  3.515 1.585 4.405 1.745 ;
        RECT  3.745 0.810 4.005 1.070 ;
        RECT  3.075 2.095 3.965 2.255 ;
        RECT  2.295 0.470 3.875 0.630 ;
        RECT  3.415 1.355 3.515 1.745 ;
        RECT  3.255 0.810 3.415 1.745 ;
        RECT  2.635 0.810 3.255 0.970 ;
        RECT  2.915 1.150 3.075 2.255 ;
        RECT  2.815 1.150 2.915 1.310 ;
        RECT  2.755 2.095 2.915 2.255 ;
        RECT  2.475 0.810 2.635 1.085 ;
        RECT  1.775 0.925 2.475 1.085 ;
        RECT  2.135 0.470 2.295 0.745 ;
        RECT  0.725 0.585 2.135 0.745 ;
        RECT  1.775 2.060 2.075 2.220 ;
        RECT  1.615 0.925 1.775 2.220 ;
        RECT  1.415 2.775 1.675 3.035 ;
        RECT  1.335 2.775 1.415 2.935 ;
        RECT  1.115 1.035 1.365 1.295 ;
        RECT  1.175 2.195 1.335 2.935 ;
        RECT  1.115 2.195 1.175 2.355 ;
        RECT  1.105 1.035 1.115 2.355 ;
        RECT  0.955 1.135 1.105 2.355 ;
        RECT  0.565 0.585 0.725 2.355 ;
        RECT  0.125 0.910 0.565 1.170 ;
        RECT  0.385 2.195 0.565 2.355 ;
        RECT  0.125 2.195 0.385 2.455 ;
    END
END SDFFHQX8

MACRO SDFFHQX4
    CLASS CORE ;
    FOREIGN SDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.085 1.235 5.395 1.990 ;
        END
        ANTENNAGATEAREA     0.1443 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.575 2.225 1.835 ;
        RECT  1.965 1.290 2.175 1.835 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.500 1.515 14.595 2.585 ;
        RECT  14.240 0.595 14.500 3.060 ;
        END
        ANTENNADIFFAREA     0.8132 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.545 2.705 1.915 ;
        RECT  2.545 1.290 2.635 1.915 ;
        RECT  2.450 1.290 2.545 1.705 ;
        RECT  2.425 1.290 2.450 1.580 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.455 0.385 2.015 ;
        END
        ANTENNAGATEAREA     0.3731 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.010 -0.250 15.180 0.250 ;
        RECT  14.750 -0.250 15.010 1.095 ;
        RECT  13.990 -0.250 14.750 0.250 ;
        RECT  13.730 -0.250 13.990 0.755 ;
        RECT  13.005 -0.250 13.730 0.250 ;
        RECT  12.745 -0.250 13.005 0.950 ;
        RECT  10.230 -0.250 12.745 0.250 ;
        RECT  9.970 -0.250 10.230 0.405 ;
        RECT  9.290 -0.250 9.970 0.250 ;
        RECT  9.030 -0.250 9.290 0.405 ;
        RECT  8.185 -0.250 9.030 0.250 ;
        RECT  7.925 -0.250 8.185 0.405 ;
        RECT  6.545 -0.250 7.925 0.250 ;
        RECT  6.385 -0.250 6.545 1.070 ;
        RECT  4.985 -0.250 6.385 0.250 ;
        RECT  6.195 0.810 6.385 1.070 ;
        RECT  4.725 -0.250 4.985 0.625 ;
        RECT  1.955 -0.250 4.725 0.250 ;
        RECT  1.695 -0.250 1.955 0.405 ;
        RECT  0.815 -0.250 1.695 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.035 3.440 15.180 3.940 ;
        RECT  14.775 2.275 15.035 3.940 ;
        RECT  13.990 3.440 14.775 3.940 ;
        RECT  13.390 2.955 13.990 3.940 ;
        RECT  10.285 3.440 13.390 3.940 ;
        RECT  10.025 3.285 10.285 3.940 ;
        RECT  9.195 3.440 10.025 3.940 ;
        RECT  8.935 3.285 9.195 3.940 ;
        RECT  7.605 3.440 8.935 3.940 ;
        RECT  7.345 3.285 7.605 3.940 ;
        RECT  6.135 3.440 7.345 3.940 ;
        RECT  5.875 3.285 6.135 3.940 ;
        RECT  5.335 3.440 5.875 3.940 ;
        RECT  5.075 3.285 5.335 3.940 ;
        RECT  3.415 3.440 5.075 3.940 ;
        RECT  2.475 3.115 3.415 3.940 ;
        RECT  0.725 3.440 2.475 3.940 ;
        RECT  0.125 2.805 0.725 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.875 1.510 13.975 1.770 ;
        RECT  13.715 1.510 13.875 2.730 ;
        RECT  12.555 2.570 13.715 2.730 ;
        RECT  13.465 1.035 13.515 1.295 ;
        RECT  13.465 2.040 13.505 2.300 ;
        RECT  13.305 1.035 13.465 2.300 ;
        RECT  13.255 1.035 13.305 1.295 ;
        RECT  12.990 1.540 13.305 1.700 ;
        RECT  13.245 2.040 13.305 2.300 ;
        RECT  12.730 1.490 12.990 1.750 ;
        RECT  12.550 2.065 12.785 2.325 ;
        RECT  12.115 2.505 12.555 2.765 ;
        RECT  12.390 0.470 12.550 2.325 ;
        RECT  12.215 2.960 12.475 3.220 ;
        RECT  10.570 0.470 12.390 0.630 ;
        RECT  10.625 3.060 12.215 3.220 ;
        RECT  12.050 1.150 12.210 1.530 ;
        RECT  11.955 2.165 12.115 2.765 ;
        RECT  11.250 1.150 12.050 1.310 ;
        RECT  11.250 2.165 11.955 2.325 ;
        RECT  10.910 0.810 11.860 0.970 ;
        RECT  11.445 2.505 11.705 2.765 ;
        RECT  10.685 2.605 11.445 2.765 ;
        RECT  11.195 1.150 11.250 2.325 ;
        RECT  11.090 1.150 11.195 2.425 ;
        RECT  10.935 2.165 11.090 2.425 ;
        RECT  10.750 0.810 10.910 1.085 ;
        RECT  10.740 0.925 10.750 1.085 ;
        RECT  10.480 0.925 10.740 1.185 ;
        RECT  10.425 2.505 10.685 2.765 ;
        RECT  10.465 2.945 10.625 3.220 ;
        RECT  10.410 0.470 10.570 0.745 ;
        RECT  9.915 0.925 10.480 1.085 ;
        RECT  8.825 2.945 10.465 3.105 ;
        RECT  9.745 2.605 10.425 2.765 ;
        RECT  6.885 0.585 10.410 0.745 ;
        RECT  9.755 0.925 9.915 2.170 ;
        RECT  9.570 0.925 9.755 1.185 ;
        RECT  9.745 2.010 9.755 2.170 ;
        RECT  9.485 2.010 9.745 2.765 ;
        RECT  9.380 1.515 9.575 1.775 ;
        RECT  8.965 2.010 9.485 2.170 ;
        RECT  9.220 0.955 9.380 1.775 ;
        RECT  8.255 0.955 9.220 1.115 ;
        RECT  8.805 1.535 8.965 2.170 ;
        RECT  8.565 2.845 8.825 3.105 ;
        RECT  8.705 1.535 8.805 1.795 ;
        RECT  6.285 2.945 8.565 3.105 ;
        RECT  8.255 2.405 8.455 2.665 ;
        RECT  8.095 0.955 8.255 2.710 ;
        RECT  7.065 0.955 8.095 1.115 ;
        RECT  6.755 2.550 8.095 2.710 ;
        RECT  7.170 1.905 7.430 2.165 ;
        RECT  6.885 1.905 7.170 2.065 ;
        RECT  6.725 0.585 6.885 2.065 ;
        RECT  6.495 2.500 6.755 2.760 ;
        RECT  5.945 1.250 6.725 1.410 ;
        RECT  6.285 1.590 6.385 1.850 ;
        RECT  6.125 1.590 6.285 3.105 ;
        RECT  5.335 0.470 6.205 0.630 ;
        RECT  4.675 2.945 6.125 3.105 ;
        RECT  5.735 0.865 5.945 1.410 ;
        RECT  5.575 0.865 5.735 2.765 ;
        RECT  5.475 2.215 5.575 2.765 ;
        RECT  1.675 2.435 5.475 2.595 ;
        RECT  5.175 0.470 5.335 0.970 ;
        RECT  4.905 0.810 5.175 0.970 ;
        RECT  4.745 0.810 4.905 2.255 ;
        RECT  4.020 0.810 4.745 0.970 ;
        RECT  4.215 2.095 4.745 2.255 ;
        RECT  4.515 2.775 4.675 3.105 ;
        RECT  4.405 1.585 4.565 1.845 ;
        RECT  1.675 2.775 4.515 2.935 ;
        RECT  3.515 1.585 4.405 1.745 ;
        RECT  3.860 0.810 4.020 1.110 ;
        RECT  3.075 2.095 3.965 2.255 ;
        RECT  2.295 0.470 3.875 0.630 ;
        RECT  3.760 0.850 3.860 1.110 ;
        RECT  3.415 1.355 3.515 1.745 ;
        RECT  3.255 0.810 3.415 1.745 ;
        RECT  2.635 0.810 3.255 0.970 ;
        RECT  2.915 1.150 3.075 2.255 ;
        RECT  2.815 1.150 2.915 1.310 ;
        RECT  2.755 2.095 2.915 2.255 ;
        RECT  2.475 0.810 2.635 1.085 ;
        RECT  1.775 0.925 2.475 1.085 ;
        RECT  2.135 0.470 2.295 0.745 ;
        RECT  0.775 0.585 2.135 0.745 ;
        RECT  1.775 2.060 2.075 2.220 ;
        RECT  1.615 0.925 1.775 2.220 ;
        RECT  1.415 2.775 1.675 3.035 ;
        RECT  1.115 2.775 1.415 2.935 ;
        RECT  1.315 0.965 1.365 1.225 ;
        RECT  1.115 0.965 1.315 1.295 ;
        RECT  1.105 0.965 1.115 2.935 ;
        RECT  0.955 1.135 1.105 2.935 ;
        RECT  0.615 0.585 0.775 2.385 ;
        RECT  0.125 0.900 0.615 1.160 ;
        RECT  0.385 2.225 0.615 2.385 ;
        RECT  0.125 2.225 0.385 2.485 ;
    END
END SDFFHQX4

MACRO SDFFHQX2
    CLASS CORE ;
    FOREIGN SDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.535 1.465 4.935 1.990 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.520 2.055 2.780 ;
        RECT  1.505 2.520 1.715 2.810 ;
        END
        ANTENNAGATEAREA     0.1729 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.825 0.695 11.835 2.995 ;
        RECT  11.565 0.600 11.825 3.055 ;
        END
        ANTENNADIFFAREA     0.7276 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.265 2.595 1.580 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.455 0.335 2.015 ;
        END
        ANTENNAGATEAREA     0.2353 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.315 -0.250 11.960 0.250 ;
        RECT  11.055 -0.250 11.315 1.095 ;
        RECT  10.025 -0.250 11.055 0.250 ;
        RECT  9.765 -0.250 10.025 1.045 ;
        RECT  7.975 -0.250 9.765 0.250 ;
        RECT  7.715 -0.250 7.975 0.405 ;
        RECT  6.835 -0.250 7.715 0.250 ;
        RECT  6.575 -0.250 6.835 0.405 ;
        RECT  4.665 -0.250 6.575 0.250 ;
        RECT  4.405 -0.250 4.665 0.790 ;
        RECT  2.495 -0.250 4.405 0.250 ;
        RECT  2.235 -0.250 2.495 0.405 ;
        RECT  0.335 -0.250 2.235 0.250 ;
        RECT  0.175 -0.250 0.335 0.690 ;
        RECT  0.000 -0.250 0.175 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.315 3.440 11.960 3.940 ;
        RECT  10.715 2.955 11.315 3.940 ;
        RECT  8.355 3.440 10.715 3.940 ;
        RECT  8.095 3.285 8.355 3.940 ;
        RECT  7.405 3.440 8.095 3.940 ;
        RECT  7.145 3.285 7.405 3.940 ;
        RECT  5.905 3.440 7.145 3.940 ;
        RECT  5.645 3.285 5.905 3.940 ;
        RECT  4.855 3.440 5.645 3.940 ;
        RECT  4.595 3.285 4.855 3.940 ;
        RECT  2.345 3.440 4.595 3.940 ;
        RECT  2.185 3.065 2.345 3.940 ;
        RECT  0.675 3.440 2.185 3.940 ;
        RECT  0.415 2.780 0.675 3.940 ;
        RECT  0.000 3.440 0.415 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.045 1.510 11.205 2.575 ;
        RECT  10.945 1.510 11.045 1.770 ;
        RECT  9.885 2.415 11.045 2.575 ;
        RECT  10.720 1.955 10.825 2.215 ;
        RECT  10.720 1.035 10.725 1.295 ;
        RECT  10.560 1.035 10.720 2.215 ;
        RECT  10.465 1.035 10.560 1.675 ;
        RECT  10.375 1.415 10.465 1.675 ;
        RECT  9.935 1.225 10.095 2.045 ;
        RECT  9.380 1.225 9.935 1.385 ;
        RECT  9.715 2.315 9.885 2.575 ;
        RECT  9.555 1.615 9.715 2.575 ;
        RECT  9.040 1.615 9.555 1.775 ;
        RECT  8.865 2.415 9.555 2.575 ;
        RECT  9.110 2.775 9.545 3.035 ;
        RECT  9.220 0.470 9.380 1.385 ;
        RECT  9.115 1.955 9.375 2.215 ;
        RECT  8.320 0.470 9.220 0.630 ;
        RECT  8.565 1.955 9.115 2.115 ;
        RECT  8.945 2.775 9.110 3.105 ;
        RECT  8.880 0.960 9.040 1.775 ;
        RECT  7.035 2.945 8.945 3.105 ;
        RECT  8.780 0.960 8.880 1.220 ;
        RECT  8.605 2.315 8.865 2.575 ;
        RECT  8.530 1.035 8.565 2.115 ;
        RECT  8.405 0.935 8.530 2.115 ;
        RECT  8.270 0.935 8.405 1.195 ;
        RECT  7.955 1.955 8.405 2.115 ;
        RECT  8.160 0.470 8.320 0.745 ;
        RECT  8.175 1.405 8.225 1.665 ;
        RECT  8.090 1.405 8.175 1.675 ;
        RECT  6.115 0.585 8.160 0.745 ;
        RECT  7.930 1.025 8.090 1.675 ;
        RECT  7.795 1.955 7.955 2.765 ;
        RECT  7.235 1.025 7.930 1.185 ;
        RECT  7.695 1.960 7.795 2.765 ;
        RECT  7.345 1.960 7.695 2.120 ;
        RECT  7.185 1.465 7.345 2.120 ;
        RECT  6.975 0.925 7.235 1.185 ;
        RECT  7.085 1.465 7.185 1.725 ;
        RECT  6.775 2.805 7.035 3.105 ;
        RECT  6.515 1.025 6.975 1.185 ;
        RECT  2.685 2.945 6.775 3.105 ;
        RECT  6.515 2.025 6.615 2.625 ;
        RECT  6.355 1.025 6.515 2.625 ;
        RECT  5.695 1.150 6.355 1.310 ;
        RECT  5.955 0.585 6.115 0.970 ;
        RECT  5.445 0.810 5.955 0.970 ;
        RECT  5.445 1.645 5.840 1.905 ;
        RECT  5.005 0.470 5.660 0.630 ;
        RECT  5.395 0.810 5.445 2.300 ;
        RECT  5.285 0.810 5.395 2.765 ;
        RECT  5.185 0.995 5.285 1.255 ;
        RECT  5.135 2.140 5.285 2.765 ;
        RECT  3.025 2.605 5.135 2.765 ;
        RECT  4.845 0.470 5.005 1.200 ;
        RECT  4.355 1.040 4.845 1.200 ;
        RECT  4.195 1.040 4.355 2.375 ;
        RECT  3.840 0.430 4.225 0.590 ;
        RECT  3.595 1.040 4.195 1.300 ;
        RECT  3.665 2.215 4.195 2.375 ;
        RECT  3.855 1.650 4.015 2.030 ;
        RECT  3.415 1.650 3.855 1.810 ;
        RECT  3.680 0.430 3.840 0.745 ;
        RECT  2.035 0.585 3.680 0.745 ;
        RECT  3.255 0.925 3.415 1.810 ;
        RECT  3.205 2.045 3.365 2.400 ;
        RECT  1.695 0.925 3.255 1.085 ;
        RECT  3.075 2.045 3.205 2.205 ;
        RECT  2.915 1.265 3.075 2.205 ;
        RECT  2.865 2.385 3.025 2.765 ;
        RECT  2.775 1.265 2.915 1.425 ;
        RECT  2.735 2.385 2.865 2.545 ;
        RECT  2.575 1.815 2.735 2.545 ;
        RECT  2.525 2.725 2.685 3.105 ;
        RECT  1.695 1.815 2.575 1.975 ;
        RECT  2.395 2.725 2.525 2.885 ;
        RECT  2.235 2.180 2.395 2.885 ;
        RECT  1.355 2.180 2.235 2.340 ;
        RECT  1.875 0.470 2.035 0.745 ;
        RECT  0.675 0.470 1.875 0.630 ;
        RECT  1.015 3.025 1.825 3.185 ;
        RECT  1.535 0.810 1.695 1.085 ;
        RECT  1.535 1.695 1.695 1.975 ;
        RECT  1.015 0.810 1.535 0.970 ;
        RECT  1.195 1.150 1.355 2.340 ;
        RECT  0.855 0.810 1.015 3.185 ;
        RECT  0.515 0.470 0.675 2.360 ;
        RECT  0.125 1.015 0.515 1.275 ;
        RECT  0.385 2.200 0.515 2.360 ;
        RECT  0.125 2.200 0.385 2.460 ;
    END
END SDFFHQX2

MACRO SDFFHQX1
    CLASS CORE ;
    FOREIGN SDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.725 1.700 4.935 1.990 ;
        RECT  4.495 1.765 4.725 1.925 ;
        RECT  4.335 1.470 4.495 1.925 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.520 2.055 2.780 ;
        RECT  1.505 2.520 1.715 2.810 ;
        END
        ANTENNAGATEAREA     0.1222 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.890 1.105 10.915 1.990 ;
        RECT  10.865 0.940 10.890 1.990 ;
        RECT  10.705 0.940 10.865 2.215 ;
        RECT  10.435 0.840 10.705 1.100 ;
        RECT  10.605 1.955 10.705 2.215 ;
        END
        ANTENNADIFFAREA     0.3876 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.265 2.625 1.580 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.475 0.335 2.020 ;
        END
        ANTENNAGATEAREA     0.1456 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.715 -0.250 11.040 0.250 ;
        RECT  10.355 -0.250 10.715 0.405 ;
        RECT  9.505 -0.250 10.355 0.250 ;
        RECT  9.245 -0.250 9.505 0.405 ;
        RECT  7.705 -0.250 9.245 0.250 ;
        RECT  7.445 -0.250 7.705 0.405 ;
        RECT  6.455 -0.250 7.445 0.250 ;
        RECT  6.195 -0.250 6.455 0.405 ;
        RECT  4.450 -0.250 6.195 0.250 ;
        RECT  4.290 -0.250 4.450 0.745 ;
        RECT  2.525 -0.250 4.290 0.250 ;
        RECT  2.265 -0.250 2.525 0.405 ;
        RECT  0.335 -0.250 2.265 0.250 ;
        RECT  0.175 -0.250 0.335 0.785 ;
        RECT  0.000 -0.250 0.175 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.325 3.440 11.040 3.940 ;
        RECT  10.065 2.870 10.325 3.940 ;
        RECT  7.945 3.440 10.065 3.940 ;
        RECT  6.885 3.285 7.945 3.940 ;
        RECT  5.385 3.440 6.885 3.940 ;
        RECT  5.125 3.285 5.385 3.940 ;
        RECT  4.435 3.440 5.125 3.940 ;
        RECT  4.175 3.285 4.435 3.940 ;
        RECT  2.085 3.440 4.175 3.940 ;
        RECT  1.925 2.990 2.085 3.940 ;
        RECT  0.675 3.440 1.925 3.940 ;
        RECT  0.415 2.735 0.675 3.940 ;
        RECT  0.000 3.440 0.415 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.795 3.025 10.895 3.185 ;
        RECT  10.635 2.430 10.795 3.185 ;
        RECT  10.095 2.430 10.635 2.590 ;
        RECT  10.095 1.405 10.155 1.665 ;
        RECT  9.935 0.905 10.095 2.590 ;
        RECT  9.895 0.905 9.935 1.665 ;
        RECT  9.890 0.905 9.895 1.615 ;
        RECT  9.835 0.905 9.890 1.165 ;
        RECT  9.465 1.225 9.625 2.015 ;
        RECT  9.375 2.990 9.520 3.150 ;
        RECT  9.375 2.245 9.475 2.505 ;
        RECT  9.105 1.225 9.465 1.385 ;
        RECT  9.255 2.245 9.375 3.150 ;
        RECT  9.215 1.565 9.255 3.150 ;
        RECT  9.095 1.565 9.215 2.725 ;
        RECT  8.945 0.635 9.105 1.385 ;
        RECT  8.765 1.565 9.095 1.725 ;
        RECT  8.455 2.565 9.095 2.725 ;
        RECT  8.600 0.635 8.945 0.795 ;
        RECT  8.755 1.905 8.915 2.385 ;
        RECT  8.535 2.905 8.795 3.165 ;
        RECT  8.605 0.980 8.765 1.725 ;
        RECT  8.295 1.905 8.755 2.065 ;
        RECT  8.505 0.980 8.605 1.240 ;
        RECT  8.340 0.535 8.600 0.795 ;
        RECT  6.455 2.905 8.535 3.065 ;
        RECT  8.295 2.245 8.455 2.725 ;
        RECT  7.165 0.635 8.340 0.795 ;
        RECT  8.135 1.025 8.295 2.065 ;
        RECT  8.195 2.245 8.295 2.505 ;
        RECT  7.995 1.025 8.135 1.285 ;
        RECT  7.545 1.905 8.135 2.065 ;
        RECT  7.695 1.465 7.955 1.725 ;
        RECT  7.515 1.465 7.695 1.625 ;
        RECT  7.285 1.905 7.545 2.425 ;
        RECT  7.355 1.150 7.515 1.625 ;
        RECT  6.965 1.150 7.355 1.310 ;
        RECT  6.990 1.905 7.285 2.065 ;
        RECT  6.905 0.535 7.165 0.795 ;
        RECT  6.830 1.515 6.990 2.065 ;
        RECT  6.705 1.035 6.965 1.310 ;
        RECT  6.195 0.635 6.905 0.795 ;
        RECT  6.595 1.515 6.830 1.675 ;
        RECT  5.935 1.150 6.705 1.310 ;
        RECT  6.405 2.785 6.455 3.065 ;
        RECT  6.195 2.785 6.405 3.105 ;
        RECT  6.205 2.275 6.255 2.535 ;
        RECT  5.995 2.155 6.205 2.535 ;
        RECT  6.035 0.635 6.195 0.970 ;
        RECT  2.425 2.945 6.195 3.105 ;
        RECT  5.275 0.810 6.035 0.970 ;
        RECT  5.935 2.155 5.995 2.315 ;
        RECT  5.775 1.150 5.935 2.315 ;
        RECT  5.485 1.150 5.775 1.310 ;
        RECT  5.275 1.715 5.595 1.975 ;
        RECT  4.790 0.470 5.340 0.630 ;
        RECT  5.115 0.810 5.275 2.330 ;
        RECT  4.975 1.035 5.115 1.295 ;
        RECT  5.025 2.170 5.115 2.330 ;
        RECT  4.925 2.170 5.025 2.430 ;
        RECT  4.765 2.170 4.925 2.765 ;
        RECT  4.630 0.470 4.790 1.085 ;
        RECT  2.765 2.605 4.765 2.765 ;
        RECT  4.155 0.925 4.630 1.085 ;
        RECT  3.995 0.925 4.155 2.325 ;
        RECT  3.850 0.470 4.110 0.745 ;
        RECT  3.655 1.035 3.995 1.295 ;
        RECT  3.665 2.165 3.995 2.325 ;
        RECT  2.095 0.585 3.850 0.745 ;
        RECT  3.445 1.825 3.815 1.985 ;
        RECT  3.405 2.165 3.665 2.425 ;
        RECT  3.285 0.925 3.445 1.985 ;
        RECT  1.720 0.925 3.285 1.085 ;
        RECT  2.945 1.265 3.105 2.425 ;
        RECT  2.805 1.265 2.945 1.425 ;
        RECT  2.605 1.815 2.765 2.765 ;
        RECT  1.725 1.815 2.605 1.975 ;
        RECT  2.265 2.180 2.425 3.105 ;
        RECT  1.355 2.180 2.265 2.340 ;
        RECT  1.935 0.470 2.095 0.745 ;
        RECT  0.675 0.470 1.935 0.630 ;
        RECT  1.565 1.715 1.725 1.975 ;
        RECT  1.560 0.810 1.720 1.085 ;
        RECT  1.015 3.000 1.565 3.160 ;
        RECT  1.015 0.810 1.560 0.970 ;
        RECT  1.195 1.150 1.355 2.340 ;
        RECT  0.855 0.810 1.015 3.160 ;
        RECT  0.515 0.470 0.675 2.360 ;
        RECT  0.125 1.035 0.515 1.295 ;
        RECT  0.385 2.200 0.515 2.360 ;
        RECT  0.125 2.200 0.385 2.460 ;
    END
END SDFFHQX1

MACRO MDFFHQX8
    CLASS CORE ;
    FOREIGN MDFFHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.905 1.680 3.220 1.990 ;
        RECT  2.745 1.485 2.905 1.990 ;
        RECT  2.410 1.485 2.745 1.645 ;
        RECT  2.250 0.585 2.410 1.645 ;
        RECT  1.595 0.585 2.250 0.745 ;
        RECT  1.335 0.430 1.595 0.745 ;
        END
        ANTENNAGATEAREA     0.6513 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.760 0.695 17.815 2.585 ;
        RECT  17.500 0.600 17.760 3.050 ;
        RECT  16.740 1.195 17.500 1.990 ;
        RECT  16.480 0.600 16.740 3.050 ;
        END
        ANTENNADIFFAREA     1.5960 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.570 1.165 0.945 1.710 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.060 1.200 5.395 1.725 ;
        END
        ANTENNAGATEAREA     0.2730 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.160 6.920 1.420 ;
        RECT  6.565 1.160 6.775 1.580 ;
        RECT  5.980 1.160 6.565 1.420 ;
        END
        ANTENNAGATEAREA     0.4238 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.270 -0.250 18.400 0.250 ;
        RECT  18.010 -0.250 18.270 1.210 ;
        RECT  17.250 -0.250 18.010 0.250 ;
        RECT  16.990 -0.250 17.250 0.965 ;
        RECT  16.200 -0.250 16.990 0.250 ;
        RECT  15.940 -0.250 16.200 0.405 ;
        RECT  15.400 -0.250 15.940 0.250 ;
        RECT  15.140 -0.250 15.400 0.405 ;
        RECT  12.600 -0.250 15.140 0.250 ;
        RECT  12.340 -0.250 12.600 0.785 ;
        RECT  11.520 -0.250 12.340 0.250 ;
        RECT  11.260 -0.250 11.520 0.865 ;
        RECT  10.325 -0.250 11.260 0.250 ;
        RECT  10.065 -0.250 10.325 0.405 ;
        RECT  8.560 -0.250 10.065 0.250 ;
        RECT  8.300 -0.250 8.560 0.405 ;
        RECT  7.160 -0.250 8.300 0.250 ;
        RECT  6.900 -0.250 7.160 0.405 ;
        RECT  6.080 -0.250 6.900 0.250 ;
        RECT  5.820 -0.250 6.080 0.405 ;
        RECT  5.030 -0.250 5.820 0.250 ;
        RECT  4.770 -0.250 5.030 0.795 ;
        RECT  3.470 -0.250 4.770 0.250 ;
        RECT  3.210 -0.250 3.470 0.895 ;
        RECT  2.410 -0.250 3.210 0.250 ;
        RECT  2.150 -0.250 2.410 0.405 ;
        RECT  1.020 -0.250 2.150 0.250 ;
        RECT  0.760 -0.250 1.020 0.405 ;
        RECT  0.000 -0.250 0.760 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.270 3.440 18.400 3.940 ;
        RECT  18.010 2.060 18.270 3.940 ;
        RECT  17.250 3.440 18.010 3.940 ;
        RECT  16.990 2.255 17.250 3.940 ;
        RECT  16.225 3.440 16.990 3.940 ;
        RECT  15.965 2.595 16.225 3.940 ;
        RECT  15.350 3.440 15.965 3.940 ;
        RECT  15.090 2.475 15.350 3.940 ;
        RECT  12.650 3.440 15.090 3.940 ;
        RECT  12.390 3.285 12.650 3.940 ;
        RECT  11.570 3.440 12.390 3.940 ;
        RECT  11.310 3.285 11.570 3.940 ;
        RECT  10.300 3.440 11.310 3.940 ;
        RECT  10.040 2.890 10.300 3.940 ;
        RECT  8.590 3.440 10.040 3.940 ;
        RECT  8.330 3.285 8.590 3.940 ;
        RECT  7.500 3.440 8.330 3.940 ;
        RECT  7.240 3.285 7.500 3.940 ;
        RECT  5.550 3.440 7.240 3.940 ;
        RECT  5.290 3.285 5.550 3.940 ;
        RECT  4.100 3.440 5.290 3.940 ;
        RECT  3.840 2.895 4.100 3.940 ;
        RECT  3.000 3.440 3.840 3.940 ;
        RECT  2.740 2.895 3.000 3.940 ;
        RECT  1.440 3.440 2.740 3.940 ;
        RECT  1.180 3.285 1.440 3.940 ;
        RECT  0.000 3.440 1.180 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.195 1.490 16.295 1.750 ;
        RECT  16.035 0.585 16.195 1.750 ;
        RECT  14.500 0.585 16.035 0.745 ;
        RECT  15.730 1.035 15.830 1.295 ;
        RECT  15.730 1.955 15.830 2.215 ;
        RECT  15.570 1.035 15.730 2.215 ;
        RECT  14.940 1.555 15.570 1.820 ;
        RECT  14.600 0.955 14.760 3.100 ;
        RECT  14.490 0.955 14.600 1.215 ;
        RECT  10.740 2.940 14.600 3.100 ;
        RECT  14.310 0.515 14.500 0.775 ;
        RECT  14.310 1.955 14.420 2.215 ;
        RECT  14.260 0.515 14.310 2.215 ;
        RECT  14.240 0.515 14.260 2.115 ;
        RECT  14.150 0.585 14.240 2.115 ;
        RECT  13.510 0.585 14.150 0.745 ;
        RECT  13.560 1.955 14.150 2.115 ;
        RECT  13.810 2.465 14.070 2.725 ;
        RECT  13.810 1.035 13.970 1.605 ;
        RECT  13.005 1.445 13.810 1.605 ;
        RECT  13.050 2.565 13.810 2.725 ;
        RECT  13.400 1.955 13.560 2.380 ;
        RECT  13.250 0.585 13.510 1.265 ;
        RECT  13.300 2.120 13.400 2.380 ;
        RECT  13.000 2.125 13.050 2.725 ;
        RECT  13.000 1.035 13.005 1.605 ;
        RECT  12.840 1.035 13.000 2.725 ;
        RECT  12.060 1.035 12.840 1.295 ;
        RECT  12.790 2.125 12.840 2.725 ;
        RECT  12.110 2.565 12.790 2.725 ;
        RECT  11.420 1.585 12.285 1.845 ;
        RECT  11.850 2.125 12.110 2.725 ;
        RECT  11.800 0.690 12.060 1.295 ;
        RECT  11.340 2.470 11.850 2.630 ;
        RECT  11.260 1.135 11.420 2.180 ;
        RECT  11.080 2.420 11.340 2.680 ;
        RECT  10.780 1.135 11.260 1.295 ;
        RECT  10.660 2.020 11.260 2.180 ;
        RECT  10.720 0.535 10.980 0.795 ;
        RECT  10.520 1.035 10.780 1.295 ;
        RECT  10.580 2.550 10.740 3.100 ;
        RECT  9.780 0.635 10.720 0.795 ;
        RECT  10.400 2.020 10.660 2.280 ;
        RECT  10.345 1.475 10.605 1.735 ;
        RECT  9.845 2.550 10.580 2.710 ;
        RECT  9.440 1.035 10.520 1.195 ;
        RECT  9.440 2.020 10.400 2.180 ;
        RECT  9.000 1.475 10.345 1.635 ;
        RECT  9.685 2.550 9.845 2.765 ;
        RECT  9.620 0.430 9.780 0.795 ;
        RECT  9.000 2.605 9.685 2.765 ;
        RECT  9.000 0.430 9.620 0.590 ;
        RECT  9.010 2.945 9.610 3.215 ;
        RECT  9.280 0.770 9.440 1.195 ;
        RECT  9.230 2.020 9.440 2.420 ;
        RECT  9.180 0.770 9.280 1.030 ;
        RECT  9.180 2.160 9.230 2.420 ;
        RECT  4.460 2.945 9.010 3.105 ;
        RECT  8.840 0.430 9.000 0.745 ;
        RECT  8.840 1.245 9.000 2.765 ;
        RECT  8.290 0.585 8.840 0.745 ;
        RECT  8.760 1.245 8.840 1.405 ;
        RECT  5.735 2.605 8.840 2.765 ;
        RECT  8.500 1.145 8.760 1.405 ;
        RECT  8.290 1.610 8.660 1.885 ;
        RECT  8.130 0.585 8.290 2.285 ;
        RECT  7.730 0.885 8.130 1.145 ;
        RECT  8.050 2.125 8.130 2.285 ;
        RECT  7.790 2.125 8.050 2.385 ;
        RECT  7.525 1.650 7.880 1.935 ;
        RECT  6.090 2.225 7.790 2.385 ;
        RECT  7.365 0.710 7.525 1.935 ;
        RECT  6.620 0.710 7.365 0.870 ;
        RECT  6.300 1.775 7.365 1.935 ;
        RECT  6.360 0.610 6.620 0.870 ;
        RECT  6.040 1.775 6.300 2.040 ;
        RECT  5.575 0.710 5.735 2.765 ;
        RECT  5.540 0.710 5.575 0.870 ;
        RECT  5.280 0.610 5.540 0.870 ;
        RECT  4.800 1.955 5.010 2.555 ;
        RECT  4.750 1.610 4.800 2.555 ;
        RECT  4.640 1.610 4.750 2.120 ;
        RECT  4.440 1.610 4.640 1.770 ;
        RECT  4.440 0.495 4.490 0.755 ;
        RECT  4.300 1.950 4.460 3.105 ;
        RECT  4.280 0.495 4.440 1.770 ;
        RECT  4.195 1.950 4.300 2.670 ;
        RECT  4.230 0.495 4.280 0.755 ;
        RECT  4.090 1.950 4.195 2.110 ;
        RECT  2.475 2.510 4.195 2.670 ;
        RECT  4.050 0.935 4.090 2.110 ;
        RECT  3.930 0.495 4.050 2.110 ;
        RECT  3.720 0.495 3.930 1.095 ;
        RECT  3.590 1.275 3.750 2.330 ;
        RECT  3.510 1.275 3.590 1.495 ;
        RECT  2.565 2.170 3.590 2.330 ;
        RECT  3.350 1.120 3.510 1.495 ;
        RECT  2.960 1.120 3.350 1.280 ;
        RECT  2.800 0.810 2.960 1.280 ;
        RECT  2.700 0.810 2.800 1.070 ;
        RECT  2.405 1.825 2.565 2.330 ;
        RECT  2.225 2.510 2.475 2.765 ;
        RECT  2.065 1.825 2.225 2.765 ;
        RECT  1.815 2.945 2.075 3.165 ;
        RECT  1.935 1.825 2.065 1.985 ;
        RECT  0.390 2.605 2.065 2.765 ;
        RECT  1.775 0.940 1.935 1.985 ;
        RECT  1.425 2.165 1.885 2.425 ;
        RECT  0.730 2.945 1.815 3.105 ;
        RECT  1.675 0.940 1.775 1.495 ;
        RECT  1.265 1.035 1.425 2.425 ;
        RECT  1.165 1.035 1.265 1.295 ;
        RECT  0.730 2.265 1.265 2.425 ;
        RECT  0.570 2.015 0.730 2.425 ;
        RECT  0.470 2.945 0.730 3.165 ;
        RECT  0.390 2.015 0.570 2.175 ;
        RECT  0.230 1.005 0.390 2.175 ;
        RECT  0.230 2.355 0.390 2.765 ;
        RECT  0.130 1.005 0.230 1.265 ;
        RECT  0.130 2.355 0.230 2.615 ;
    END
END MDFFHQX8

MACRO MDFFHQX4
    CLASS CORE ;
    FOREIGN MDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.410 3.375 1.990 ;
        RECT  2.605 1.410 2.885 1.570 ;
        RECT  2.445 0.585 2.605 1.570 ;
        RECT  1.700 0.585 2.445 0.745 ;
        RECT  1.440 0.430 1.700 0.745 ;
        END
        ANTENNAGATEAREA     0.6513 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.845 1.105 16.895 2.585 ;
        RECT  16.585 0.615 16.845 3.055 ;
        END
        ANTENNADIFFAREA     0.7980 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.415 1.220 1.675 ;
        RECT  0.585 1.290 1.045 1.725 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.125 1.230 5.440 1.835 ;
        END
        ANTENNAGATEAREA     0.2730 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.160 6.980 1.420 ;
        RECT  6.565 1.160 6.775 1.580 ;
        RECT  6.040 1.160 6.565 1.420 ;
        END
        ANTENNAGATEAREA     0.4238 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.355 -0.250 17.480 0.250 ;
        RECT  17.095 -0.250 17.355 1.115 ;
        RECT  16.305 -0.250 17.095 0.250 ;
        RECT  16.045 -0.250 16.305 0.405 ;
        RECT  15.505 -0.250 16.045 0.250 ;
        RECT  15.245 -0.250 15.505 0.405 ;
        RECT  12.705 -0.250 15.245 0.250 ;
        RECT  12.445 -0.250 12.705 0.785 ;
        RECT  11.625 -0.250 12.445 0.250 ;
        RECT  11.365 -0.250 11.625 0.865 ;
        RECT  10.430 -0.250 11.365 0.250 ;
        RECT  10.170 -0.250 10.430 0.405 ;
        RECT  8.665 -0.250 10.170 0.250 ;
        RECT  8.405 -0.250 8.665 0.405 ;
        RECT  7.265 -0.250 8.405 0.250 ;
        RECT  7.005 -0.250 7.265 0.405 ;
        RECT  6.185 -0.250 7.005 0.250 ;
        RECT  5.925 -0.250 6.185 0.405 ;
        RECT  5.135 -0.250 5.925 0.250 ;
        RECT  4.875 -0.250 5.135 0.795 ;
        RECT  3.575 -0.250 4.875 0.250 ;
        RECT  3.315 -0.250 3.575 0.845 ;
        RECT  2.515 -0.250 3.315 0.250 ;
        RECT  2.255 -0.250 2.515 0.405 ;
        RECT  1.020 -0.250 2.255 0.250 ;
        RECT  0.760 -0.250 1.020 1.110 ;
        RECT  0.000 -0.250 0.760 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.355 3.440 17.480 3.940 ;
        RECT  17.095 2.255 17.355 3.940 ;
        RECT  16.330 3.440 17.095 3.940 ;
        RECT  16.070 2.595 16.330 3.940 ;
        RECT  15.455 3.440 16.070 3.940 ;
        RECT  15.195 2.475 15.455 3.940 ;
        RECT  12.755 3.440 15.195 3.940 ;
        RECT  12.495 3.285 12.755 3.940 ;
        RECT  11.675 3.440 12.495 3.940 ;
        RECT  11.415 3.285 11.675 3.940 ;
        RECT  10.405 3.440 11.415 3.940 ;
        RECT  10.145 2.890 10.405 3.940 ;
        RECT  8.695 3.440 10.145 3.940 ;
        RECT  8.435 3.285 8.695 3.940 ;
        RECT  7.605 3.440 8.435 3.940 ;
        RECT  7.345 3.285 7.605 3.940 ;
        RECT  5.655 3.440 7.345 3.940 ;
        RECT  5.395 3.285 5.655 3.940 ;
        RECT  4.105 3.440 5.395 3.940 ;
        RECT  3.845 3.285 4.105 3.940 ;
        RECT  3.025 3.440 3.845 3.940 ;
        RECT  2.765 2.895 3.025 3.940 ;
        RECT  1.435 3.440 2.765 3.940 ;
        RECT  1.175 3.285 1.435 3.940 ;
        RECT  0.000 3.440 1.175 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.300 1.490 16.400 1.750 ;
        RECT  16.140 0.585 16.300 1.750 ;
        RECT  14.605 0.585 16.140 0.745 ;
        RECT  15.835 1.035 15.935 1.295 ;
        RECT  15.835 1.955 15.935 2.215 ;
        RECT  15.675 1.035 15.835 2.215 ;
        RECT  15.045 1.555 15.675 1.820 ;
        RECT  14.705 0.955 14.865 3.065 ;
        RECT  14.595 0.955 14.705 1.215 ;
        RECT  14.440 2.905 14.705 3.065 ;
        RECT  14.415 0.515 14.605 0.775 ;
        RECT  14.415 1.955 14.525 2.215 ;
        RECT  14.180 2.905 14.440 3.165 ;
        RECT  14.365 0.515 14.415 2.215 ;
        RECT  14.345 0.515 14.365 2.115 ;
        RECT  14.255 0.585 14.345 2.115 ;
        RECT  13.615 0.585 14.255 0.745 ;
        RECT  13.665 1.955 14.255 2.115 ;
        RECT  10.845 2.905 14.180 3.065 ;
        RECT  13.915 2.465 14.175 2.725 ;
        RECT  13.915 1.035 14.075 1.605 ;
        RECT  13.110 1.445 13.915 1.605 ;
        RECT  13.155 2.565 13.915 2.725 ;
        RECT  13.455 1.955 13.665 2.380 ;
        RECT  13.355 0.585 13.615 1.265 ;
        RECT  13.405 2.120 13.455 2.380 ;
        RECT  13.105 2.125 13.155 2.725 ;
        RECT  13.105 1.035 13.110 1.605 ;
        RECT  12.945 1.035 13.105 2.725 ;
        RECT  12.165 1.035 12.945 1.295 ;
        RECT  12.895 2.125 12.945 2.725 ;
        RECT  12.215 2.565 12.895 2.725 ;
        RECT  11.525 1.585 12.390 1.845 ;
        RECT  11.955 2.125 12.215 2.725 ;
        RECT  11.905 0.690 12.165 1.295 ;
        RECT  11.445 2.565 11.955 2.725 ;
        RECT  11.365 1.135 11.525 2.180 ;
        RECT  11.185 2.360 11.445 2.725 ;
        RECT  10.885 1.135 11.365 1.295 ;
        RECT  10.765 2.020 11.365 2.180 ;
        RECT  10.760 0.535 11.020 0.795 ;
        RECT  10.625 1.035 10.885 1.295 ;
        RECT  10.685 2.550 10.845 3.065 ;
        RECT  10.505 2.020 10.765 2.280 ;
        RECT  9.885 0.635 10.760 0.795 ;
        RECT  9.950 2.550 10.685 2.710 ;
        RECT  9.545 1.035 10.625 1.195 ;
        RECT  10.280 1.475 10.540 1.735 ;
        RECT  9.545 2.020 10.505 2.180 ;
        RECT  9.105 1.475 10.280 1.635 ;
        RECT  9.790 2.550 9.950 2.765 ;
        RECT  9.725 0.430 9.885 0.795 ;
        RECT  9.105 2.605 9.790 2.765 ;
        RECT  9.105 0.430 9.725 0.590 ;
        RECT  9.115 2.945 9.715 3.215 ;
        RECT  9.385 0.770 9.545 1.195 ;
        RECT  9.335 2.020 9.545 2.420 ;
        RECT  9.285 0.770 9.385 1.030 ;
        RECT  9.285 2.160 9.335 2.420 ;
        RECT  4.605 2.945 9.115 3.105 ;
        RECT  8.945 0.430 9.105 0.745 ;
        RECT  8.945 1.245 9.105 2.765 ;
        RECT  8.395 0.585 8.945 0.745 ;
        RECT  8.865 1.245 8.945 1.405 ;
        RECT  5.840 2.605 8.945 2.765 ;
        RECT  8.605 1.145 8.865 1.405 ;
        RECT  8.395 1.610 8.765 1.885 ;
        RECT  8.235 0.585 8.395 2.285 ;
        RECT  7.835 0.885 8.235 1.145 ;
        RECT  8.155 2.125 8.235 2.285 ;
        RECT  7.895 2.125 8.155 2.385 ;
        RECT  7.630 1.650 7.985 1.935 ;
        RECT  6.195 2.225 7.895 2.385 ;
        RECT  7.470 0.710 7.630 1.935 ;
        RECT  6.725 0.710 7.470 0.870 ;
        RECT  6.405 1.775 7.470 1.935 ;
        RECT  6.465 0.610 6.725 0.870 ;
        RECT  6.145 1.775 6.405 2.040 ;
        RECT  5.680 0.710 5.840 2.765 ;
        RECT  5.645 0.710 5.680 0.870 ;
        RECT  5.485 0.555 5.645 0.870 ;
        RECT  5.385 0.555 5.485 0.815 ;
        RECT  4.945 2.165 5.115 2.765 ;
        RECT  4.855 1.610 4.945 2.765 ;
        RECT  4.785 1.610 4.855 2.330 ;
        RECT  4.545 1.610 4.785 1.770 ;
        RECT  4.445 1.950 4.605 3.105 ;
        RECT  4.545 0.495 4.595 0.755 ;
        RECT  4.385 0.495 4.545 1.770 ;
        RECT  4.345 1.950 4.445 2.890 ;
        RECT  4.335 0.495 4.385 0.755 ;
        RECT  4.195 1.950 4.345 2.110 ;
        RECT  2.515 2.530 4.345 2.690 ;
        RECT  4.155 0.935 4.195 2.110 ;
        RECT  4.035 0.585 4.155 2.110 ;
        RECT  3.995 0.585 4.035 1.095 ;
        RECT  3.825 0.585 3.995 0.845 ;
        RECT  3.715 1.275 3.855 2.350 ;
        RECT  3.695 1.025 3.715 2.350 ;
        RECT  3.555 1.025 3.695 1.545 ;
        RECT  2.705 2.190 3.695 2.350 ;
        RECT  3.135 1.025 3.555 1.185 ;
        RECT  2.855 0.805 3.135 1.185 ;
        RECT  2.805 0.810 2.855 1.185 ;
        RECT  2.545 1.815 2.705 2.350 ;
        RECT  2.445 1.815 2.545 2.075 ;
        RECT  2.265 2.530 2.515 2.765 ;
        RECT  2.105 1.340 2.265 2.765 ;
        RECT  1.855 2.945 2.115 3.160 ;
        RECT  2.070 1.340 2.105 1.500 ;
        RECT  0.385 2.605 2.105 2.765 ;
        RECT  1.810 0.945 2.070 1.500 ;
        RECT  1.765 2.165 1.925 2.425 ;
        RECT  0.725 2.945 1.855 3.105 ;
        RECT  1.560 2.215 1.765 2.425 ;
        RECT  1.400 0.975 1.560 2.425 ;
        RECT  1.300 0.975 1.400 1.235 ;
        RECT  0.725 2.265 1.400 2.425 ;
        RECT  0.565 1.955 0.725 2.425 ;
        RECT  0.465 2.945 0.725 3.160 ;
        RECT  0.385 1.955 0.565 2.115 ;
        RECT  0.225 0.975 0.385 2.115 ;
        RECT  0.225 2.360 0.385 2.765 ;
        RECT  0.125 0.975 0.225 1.235 ;
        RECT  0.125 2.360 0.225 2.620 ;
    END
END MDFFHQX4

MACRO MDFFHQX2
    CLASS CORE ;
    FOREIGN MDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 1.515 1.715 1.990 ;
        RECT  1.540 1.315 1.640 1.990 ;
        RECT  1.505 0.585 1.540 1.990 ;
        RECT  1.480 0.585 1.505 1.925 ;
        RECT  1.380 0.585 1.480 1.475 ;
        RECT  0.850 0.585 1.380 0.745 ;
        RECT  0.690 0.430 0.850 0.745 ;
        RECT  0.590 0.430 0.690 0.590 ;
        END
        ANTENNAGATEAREA     0.3549 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.655 0.595 10.915 3.050 ;
        END
        ANTENNADIFFAREA     0.7140 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.335 0.860 1.990 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.615 1.290 4.015 1.580 ;
        RECT  3.355 1.290 3.615 1.610 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.535 1.290 4.935 1.600 ;
        END
        ANTENNAGATEAREA     0.2327 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.375 -0.250 11.040 0.250 ;
        RECT  10.115 -0.250 10.375 0.405 ;
        RECT  9.575 -0.250 10.115 0.250 ;
        RECT  9.315 -0.250 9.575 0.405 ;
        RECT  7.455 -0.250 9.315 0.250 ;
        RECT  7.195 -0.250 7.455 0.755 ;
        RECT  5.805 -0.250 7.195 0.250 ;
        RECT  5.545 -0.250 5.805 0.405 ;
        RECT  4.200 -0.250 5.545 0.250 ;
        RECT  3.180 -0.250 4.200 0.405 ;
        RECT  1.400 -0.250 3.180 0.250 ;
        RECT  1.140 -0.250 1.400 0.405 ;
        RECT  0.000 -0.250 1.140 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.375 3.440 11.040 3.940 ;
        RECT  10.115 2.890 10.375 3.940 ;
        RECT  9.525 3.440 10.115 3.940 ;
        RECT  9.265 2.890 9.525 3.940 ;
        RECT  7.595 3.440 9.265 3.940 ;
        RECT  7.335 3.285 7.595 3.940 ;
        RECT  5.835 3.440 7.335 3.940 ;
        RECT  5.575 3.285 5.835 3.940 ;
        RECT  3.815 3.440 5.575 3.940 ;
        RECT  3.555 3.285 3.815 3.940 ;
        RECT  1.785 3.440 3.555 3.940 ;
        RECT  1.625 3.075 1.785 3.940 ;
        RECT  0.000 3.440 1.625 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.845 1.035 10.005 2.365 ;
        RECT  9.795 1.035 9.845 1.295 ;
        RECT  9.745 2.005 9.845 2.365 ;
        RECT  9.275 2.005 9.745 2.165 ;
        RECT  9.565 1.405 9.615 1.665 ;
        RECT  9.405 0.585 9.565 1.665 ;
        RECT  8.505 0.585 9.405 0.745 ;
        RECT  9.115 1.885 9.275 2.165 ;
        RECT  8.935 2.920 8.965 3.180 ;
        RECT  8.805 0.925 8.935 3.180 ;
        RECT  8.775 0.925 8.805 3.100 ;
        RECT  8.665 0.925 8.775 1.190 ;
        RECT  6.910 2.940 8.775 3.100 ;
        RECT  8.485 1.440 8.595 2.735 ;
        RECT  8.485 0.535 8.505 0.795 ;
        RECT  8.435 0.535 8.485 2.735 ;
        RECT  8.325 0.535 8.435 1.600 ;
        RECT  8.245 0.535 8.325 0.795 ;
        RECT  7.995 1.085 8.135 2.735 ;
        RECT  7.975 0.985 7.995 2.735 ;
        RECT  7.735 0.985 7.975 1.245 ;
        RECT  7.875 2.135 7.975 2.735 ;
        RECT  7.365 2.395 7.875 2.555 ;
        RECT  7.520 1.585 7.745 1.845 ;
        RECT  7.360 1.025 7.520 2.215 ;
        RECT  7.105 2.395 7.365 2.655 ;
        RECT  6.715 1.025 7.360 1.185 ;
        RECT  6.685 2.055 7.360 2.215 ;
        RECT  5.615 0.585 6.915 0.745 ;
        RECT  6.750 2.605 6.910 3.100 ;
        RECT  6.245 1.615 6.885 1.875 ;
        RECT  6.245 2.605 6.750 2.765 ;
        RECT  6.455 0.925 6.715 1.185 ;
        RECT  6.475 2.055 6.685 2.425 ;
        RECT  6.235 3.100 6.515 3.260 ;
        RECT  6.425 2.165 6.475 2.425 ;
        RECT  6.085 1.270 6.245 2.765 ;
        RECT  6.075 2.945 6.235 3.260 ;
        RECT  5.955 1.270 6.085 1.430 ;
        RECT  4.785 2.605 6.085 2.765 ;
        RECT  5.395 2.945 6.075 3.105 ;
        RECT  5.795 1.170 5.955 1.430 ;
        RECT  5.615 1.650 5.905 1.910 ;
        RECT  5.455 0.585 5.615 2.280 ;
        RECT  5.265 0.585 5.455 0.770 ;
        RECT  5.295 2.120 5.455 2.280 ;
        RECT  5.235 2.945 5.395 3.135 ;
        RECT  5.035 2.120 5.295 2.425 ;
        RECT  5.115 0.950 5.275 1.940 ;
        RECT  5.005 0.510 5.265 0.770 ;
        RECT  4.345 2.975 5.235 3.135 ;
        RECT  4.700 0.950 5.115 1.110 ;
        RECT  4.695 1.780 5.115 1.940 ;
        RECT  4.615 2.265 5.035 2.425 ;
        RECT  4.525 2.605 4.785 2.795 ;
        RECT  4.540 0.840 4.700 1.110 ;
        RECT  4.535 1.780 4.695 2.040 ;
        RECT  4.355 2.225 4.615 2.425 ;
        RECT  4.175 2.605 4.525 2.765 ;
        RECT  4.195 0.940 4.355 1.920 ;
        RECT  4.185 2.945 4.345 3.135 ;
        RECT  3.800 0.940 4.195 1.100 ;
        RECT  4.175 1.760 4.195 1.920 ;
        RECT  2.835 2.945 4.185 3.105 ;
        RECT  4.015 1.760 4.175 2.765 ;
        RECT  3.540 0.840 3.800 1.100 ;
        RECT  3.175 1.955 3.395 2.555 ;
        RECT  3.135 0.745 3.175 2.555 ;
        RECT  3.015 0.745 3.135 2.120 ;
        RECT  2.630 0.745 3.015 0.905 ;
        RECT  2.675 1.085 2.835 3.105 ;
        RECT  2.450 1.085 2.675 1.245 ;
        RECT  1.445 2.735 2.675 2.895 ;
        RECT  2.275 1.425 2.470 1.685 ;
        RECT  2.290 0.435 2.450 1.245 ;
        RECT  2.275 1.955 2.375 2.555 ;
        RECT  2.090 0.435 2.290 0.595 ;
        RECT  2.115 1.425 2.275 2.555 ;
        RECT  2.055 1.425 2.115 1.585 ;
        RECT  1.105 2.345 2.115 2.505 ;
        RECT  1.895 0.945 2.055 1.585 ;
        RECT  1.720 0.945 1.895 1.105 ;
        RECT  1.285 2.735 1.445 3.220 ;
        RECT  1.200 2.005 1.300 2.165 ;
        RECT  0.385 3.060 1.285 3.220 ;
        RECT  1.040 0.945 1.200 2.165 ;
        RECT  0.945 2.345 1.105 2.875 ;
        RECT  0.730 0.945 1.040 1.105 ;
        RECT  0.385 0.840 0.480 1.100 ;
        RECT  0.225 0.840 0.385 3.220 ;
        RECT  0.220 0.840 0.225 1.100 ;
        RECT  0.125 2.360 0.225 2.960 ;
    END
END MDFFHQX2

MACRO MDFFHQX1
    CLASS CORE ;
    FOREIGN MDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 0.470 1.795 0.905 ;
        END
        ANTENNAGATEAREA     0.2106 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.895 1.105 9.995 2.175 ;
        RECT  9.735 0.695 9.895 2.680 ;
        RECT  9.525 0.695 9.735 0.855 ;
        RECT  9.535 2.520 9.735 2.680 ;
        RECT  9.365 2.520 9.535 2.995 ;
        RECT  9.265 0.595 9.525 0.855 ;
        RECT  9.105 2.520 9.365 3.165 ;
        END
        ANTENNADIFFAREA     0.3808 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.550 1.255 1.990 ;
        RECT  0.855 1.550 1.045 1.810 ;
        END
        ANTENNAGATEAREA     0.0923 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.900 0.880 3.095 1.620 ;
        RECT  2.885 0.880 2.900 1.290 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.615 1.290 4.015 1.620 ;
        END
        ANTENNAGATEAREA     0.1300 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.985 -0.250 10.120 0.250 ;
        RECT  8.935 -0.250 8.985 0.405 ;
        RECT  8.775 -0.250 8.935 1.135 ;
        RECT  8.725 -0.250 8.775 0.405 ;
        RECT  6.830 -0.250 8.725 0.250 ;
        RECT  6.570 -0.250 6.830 0.405 ;
        RECT  5.150 -0.250 6.570 0.250 ;
        RECT  4.890 -0.250 5.150 0.405 ;
        RECT  3.200 -0.250 4.890 0.250 ;
        RECT  2.940 -0.250 3.200 0.405 ;
        RECT  1.295 -0.250 2.940 0.250 ;
        RECT  1.035 -0.250 1.295 1.295 ;
        RECT  0.000 -0.250 1.035 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.845 3.440 10.120 3.940 ;
        RECT  8.585 2.615 8.845 3.940 ;
        RECT  7.020 3.440 8.585 3.940 ;
        RECT  6.760 3.285 7.020 3.940 ;
        RECT  5.260 3.440 6.760 3.940 ;
        RECT  5.000 3.285 5.260 3.940 ;
        RECT  3.340 3.440 5.000 3.940 ;
        RECT  3.080 3.285 3.340 3.940 ;
        RECT  1.455 3.440 3.080 3.940 ;
        RECT  1.195 3.115 1.455 3.940 ;
        RECT  0.000 3.440 1.195 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.395 1.105 9.555 2.165 ;
        RECT  9.295 1.105 9.395 1.365 ;
        RECT  9.135 2.005 9.395 2.285 ;
        RECT  9.030 1.560 9.185 1.820 ;
        RECT  8.690 2.005 9.135 2.165 ;
        RECT  8.870 1.320 9.030 1.820 ;
        RECT  8.585 1.320 8.870 1.480 ;
        RECT  8.430 1.785 8.690 2.165 ;
        RECT  8.425 0.745 8.585 1.480 ;
        RECT  7.905 0.745 8.425 0.905 ;
        RECT  8.085 1.085 8.245 3.215 ;
        RECT  7.455 3.055 8.085 3.215 ;
        RECT  7.745 0.745 7.905 2.795 ;
        RECT  7.630 0.975 7.745 1.235 ;
        RECT  7.500 0.570 7.550 0.730 ;
        RECT  7.290 0.570 7.500 0.745 ;
        RECT  7.295 2.940 7.455 3.215 ;
        RECT  7.370 2.135 7.445 2.760 ;
        RECT  7.370 0.965 7.380 1.225 ;
        RECT  7.210 0.965 7.370 2.760 ;
        RECT  6.140 2.940 7.295 3.100 ;
        RECT  4.920 0.585 7.290 0.745 ;
        RECT  7.120 0.965 7.210 1.225 ;
        RECT  7.185 2.135 7.210 2.760 ;
        RECT  6.390 2.600 7.185 2.760 ;
        RECT  6.645 1.635 7.030 1.895 ;
        RECT  6.485 1.025 6.645 2.420 ;
        RECT  6.040 1.025 6.485 1.185 ;
        RECT  5.710 2.260 6.485 2.420 ;
        RECT  5.700 1.820 6.170 2.080 ;
        RECT  5.980 2.605 6.140 3.100 ;
        RECT  5.880 0.925 6.040 1.185 ;
        RECT  5.530 2.605 5.980 2.765 ;
        RECT  4.615 2.945 5.800 3.105 ;
        RECT  5.540 1.135 5.700 2.080 ;
        RECT  5.360 1.135 5.540 1.295 ;
        RECT  5.530 1.920 5.540 2.080 ;
        RECT  5.370 1.920 5.530 2.765 ;
        RECT  4.200 2.605 5.370 2.765 ;
        RECT  5.100 1.035 5.360 1.295 ;
        RECT  5.060 1.565 5.360 1.725 ;
        RECT  4.920 1.565 5.060 2.405 ;
        RECT  4.900 0.585 4.920 2.405 ;
        RECT  4.760 0.585 4.900 1.725 ;
        RECT  3.770 2.245 4.900 2.405 ;
        RECT  4.570 0.585 4.760 0.770 ;
        RECT  4.455 2.945 4.615 3.135 ;
        RECT  4.420 0.950 4.580 1.915 ;
        RECT  4.310 0.510 4.570 0.770 ;
        RECT  3.680 2.975 4.455 3.135 ;
        RECT  4.130 0.950 4.420 1.110 ;
        RECT  4.355 1.755 4.420 1.915 ;
        RECT  4.195 1.755 4.355 2.035 ;
        RECT  3.940 2.605 4.200 2.795 ;
        RECT  3.660 1.875 4.195 2.035 ;
        RECT  3.970 0.440 4.130 1.110 ;
        RECT  3.530 0.440 3.970 0.600 ;
        RECT  3.435 2.605 3.940 2.765 ;
        RECT  3.435 0.950 3.790 1.110 ;
        RECT  3.520 2.945 3.680 3.135 ;
        RECT  2.380 2.945 3.520 3.105 ;
        RECT  3.275 0.950 3.435 2.765 ;
        RECT  2.720 2.100 2.940 2.360 ;
        RECT  2.705 1.800 2.720 2.360 ;
        RECT  2.680 0.905 2.705 2.360 ;
        RECT  2.560 0.905 2.680 2.260 ;
        RECT  2.545 0.905 2.560 1.960 ;
        RECT  2.365 2.140 2.380 3.105 ;
        RECT  2.220 0.545 2.365 3.105 ;
        RECT  2.205 0.545 2.220 2.930 ;
        RECT  2.175 0.545 2.205 0.705 ;
        RECT  1.015 2.770 2.205 2.930 ;
        RECT  1.975 0.445 2.175 0.705 ;
        RECT  1.835 1.685 2.025 1.945 ;
        RECT  1.835 1.085 1.935 1.245 ;
        RECT  1.820 2.330 1.920 2.590 ;
        RECT  1.820 1.085 1.835 1.945 ;
        RECT  1.660 1.085 1.820 2.590 ;
        RECT  0.675 2.430 1.660 2.590 ;
        RECT  0.855 2.770 1.015 3.125 ;
        RECT  0.335 2.965 0.855 3.125 ;
        RECT  0.675 1.990 0.845 2.250 ;
        RECT  0.675 1.035 0.785 1.295 ;
        RECT  0.515 1.035 0.675 2.250 ;
        RECT  0.515 2.430 0.675 2.785 ;
        RECT  0.335 0.455 0.385 0.715 ;
        RECT  0.175 0.455 0.335 3.125 ;
        RECT  0.125 0.455 0.175 0.715 ;
    END
END MDFFHQX1

MACRO EDFFHQX8
    CLASS CORE ;
    FOREIGN EDFFHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.940 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.305 1.105 17.355 2.585 ;
        RECT  17.295 1.105 17.305 3.065 ;
        RECT  17.045 0.610 17.295 3.065 ;
        RECT  17.035 0.610 17.045 1.990 ;
        RECT  16.285 1.290 17.035 1.990 ;
        RECT  16.275 1.290 16.285 3.065 ;
        RECT  16.025 0.610 16.275 3.065 ;
        RECT  16.015 0.610 16.025 1.770 ;
        END
        ANTENNADIFFAREA     1.5960 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.415 3.045 1.950 ;
        RECT  2.175 1.415 2.885 1.575 ;
        RECT  2.170 1.290 2.175 1.580 ;
        RECT  1.965 1.270 2.170 1.580 ;
        RECT  1.910 1.270 1.965 1.575 ;
        END
        ANTENNAGATEAREA     0.2626 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.635 1.105 0.895 1.845 ;
        RECT  0.585 1.290 0.635 1.640 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.160 6.220 1.420 ;
        RECT  5.645 1.160 5.855 1.580 ;
        RECT  5.280 1.160 5.645 1.420 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.805 -0.250 17.940 0.250 ;
        RECT  17.545 -0.250 17.805 1.115 ;
        RECT  16.785 -0.250 17.545 0.250 ;
        RECT  16.525 -0.250 16.785 1.065 ;
        RECT  15.735 -0.250 16.525 0.250 ;
        RECT  15.475 -0.250 15.735 1.135 ;
        RECT  5.375 -0.250 15.475 0.250 ;
        RECT  5.115 -0.250 5.375 0.405 ;
        RECT  4.250 -0.250 5.115 0.250 ;
        RECT  3.990 -0.250 4.250 0.405 ;
        RECT  2.420 -0.250 3.990 0.250 ;
        RECT  2.160 -0.250 2.420 0.405 ;
        RECT  0.805 -0.250 2.160 0.250 ;
        RECT  0.545 -0.250 0.805 0.405 ;
        RECT  0.000 -0.250 0.545 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.815 3.440 17.940 3.940 ;
        RECT  17.555 2.275 17.815 3.940 ;
        RECT  16.795 3.440 17.555 3.940 ;
        RECT  16.535 2.275 16.795 3.940 ;
        RECT  15.725 3.440 16.535 3.940 ;
        RECT  15.565 2.275 15.725 3.940 ;
        RECT  14.545 3.440 15.565 3.940 ;
        RECT  14.285 3.285 14.545 3.940 ;
        RECT  11.755 3.440 14.285 3.940 ;
        RECT  11.495 3.285 11.755 3.940 ;
        RECT  10.675 3.440 11.495 3.940 ;
        RECT  10.415 3.285 10.675 3.940 ;
        RECT  9.405 3.440 10.415 3.940 ;
        RECT  9.145 2.890 9.405 3.940 ;
        RECT  7.695 3.440 9.145 3.940 ;
        RECT  7.435 3.285 7.695 3.940 ;
        RECT  6.605 3.440 7.435 3.940 ;
        RECT  6.345 3.285 6.605 3.940 ;
        RECT  4.655 3.440 6.345 3.940 ;
        RECT  4.395 3.285 4.655 3.940 ;
        RECT  2.865 3.440 4.395 3.940 ;
        RECT  2.605 3.285 2.865 3.940 ;
        RECT  1.295 3.440 2.605 3.940 ;
        RECT  1.035 3.285 1.295 3.940 ;
        RECT  0.000 3.440 1.035 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.380 1.490 15.820 1.750 ;
        RECT  15.220 1.490 15.380 2.950 ;
        RECT  14.960 0.940 15.225 1.200 ;
        RECT  14.350 2.790 15.220 2.950 ;
        RECT  14.960 2.320 15.040 2.580 ;
        RECT  14.800 0.940 14.960 2.580 ;
        RECT  14.705 0.940 14.800 1.100 ;
        RECT  14.755 1.555 14.800 2.580 ;
        RECT  14.535 1.555 14.755 1.890 ;
        RECT  14.545 0.470 14.705 1.100 ;
        RECT  10.430 0.470 14.545 0.630 ;
        RECT  14.190 0.810 14.350 2.950 ;
        RECT  11.885 0.810 14.190 0.970 ;
        RECT  13.445 2.625 14.190 2.785 ;
        RECT  13.845 1.150 14.005 2.385 ;
        RECT  11.665 1.150 13.845 1.310 ;
        RECT  12.805 2.225 13.845 2.385 ;
        RECT  12.095 3.060 13.725 3.220 ;
        RECT  13.495 1.520 13.655 2.040 ;
        RECT  11.325 1.520 13.495 1.680 ;
        RECT  13.185 2.575 13.445 2.835 ;
        RECT  12.295 2.600 13.185 2.760 ;
        RECT  12.545 2.125 12.805 2.385 ;
        RECT  11.215 2.160 12.545 2.320 ;
        RECT  12.035 2.500 12.295 2.760 ;
        RECT  11.935 2.940 12.095 3.220 ;
        RECT  9.845 2.940 11.935 3.100 ;
        RECT  11.505 0.885 11.665 1.310 ;
        RECT  10.935 0.885 11.505 1.045 ;
        RECT  11.165 1.225 11.325 1.680 ;
        RECT  10.955 2.125 11.215 2.725 ;
        RECT  10.755 1.225 11.165 1.385 ;
        RECT  10.415 1.585 10.985 1.845 ;
        RECT  10.185 2.410 10.955 2.570 ;
        RECT  10.595 0.810 10.755 1.385 ;
        RECT  10.085 0.810 10.595 0.970 ;
        RECT  10.270 0.430 10.430 0.630 ;
        RECT  10.255 1.150 10.415 2.180 ;
        RECT  9.640 0.430 10.270 0.590 ;
        RECT  8.375 1.150 10.255 1.310 ;
        RECT  9.765 2.020 10.255 2.180 ;
        RECT  9.825 0.770 10.085 0.970 ;
        RECT  9.685 2.550 9.845 3.100 ;
        RECT  7.395 0.810 9.825 0.970 ;
        RECT  9.505 2.020 9.765 2.315 ;
        RECT  8.105 2.550 9.685 2.710 ;
        RECT  9.480 0.430 9.640 0.630 ;
        RECT  9.280 1.555 9.540 1.815 ;
        RECT  8.545 2.020 9.505 2.180 ;
        RECT  5.715 0.470 9.480 0.630 ;
        RECT  8.105 1.555 9.280 1.715 ;
        RECT  8.115 2.945 8.715 3.215 ;
        RECT  8.285 2.020 8.545 2.315 ;
        RECT  3.880 2.945 8.115 3.105 ;
        RECT  7.945 1.245 8.105 2.765 ;
        RECT  7.865 1.245 7.945 1.410 ;
        RECT  4.220 2.605 7.945 2.765 ;
        RECT  7.605 1.150 7.865 1.410 ;
        RECT  7.395 1.650 7.765 1.910 ;
        RECT  7.235 0.810 7.395 2.290 ;
        RECT  6.885 0.810 7.235 1.075 ;
        RECT  7.155 2.130 7.235 2.290 ;
        RECT  6.895 2.130 7.155 2.390 ;
        RECT  6.630 1.650 6.985 1.935 ;
        RECT  5.535 2.230 6.895 2.390 ;
        RECT  6.835 0.815 6.885 1.075 ;
        RECT  6.470 0.810 6.630 1.935 ;
        RECT  5.895 0.810 6.470 0.970 ;
        RECT  5.315 1.775 6.470 1.935 ;
        RECT  5.555 0.470 5.715 0.745 ;
        RECT  5.100 0.585 5.555 0.745 ;
        RECT  5.055 1.775 5.315 2.060 ;
        RECT  4.940 0.585 5.100 1.210 ;
        RECT  4.665 1.050 4.940 1.210 ;
        RECT  4.500 0.555 4.760 0.815 ;
        RECT  4.405 1.050 4.665 1.310 ;
        RECT  4.220 0.655 4.500 0.815 ;
        RECT  4.060 0.655 4.220 2.765 ;
        RECT  3.720 0.685 3.880 3.105 ;
        RECT  3.360 0.685 3.720 0.845 ;
        RECT  3.595 2.200 3.720 2.800 ;
        RECT  2.355 2.585 3.595 2.745 ;
        RECT  3.385 1.315 3.525 1.575 ;
        RECT  3.225 1.070 3.385 2.405 ;
        RECT  3.100 0.585 3.360 0.845 ;
        RECT  2.920 1.070 3.225 1.230 ;
        RECT  2.625 2.245 3.225 2.405 ;
        RECT  2.760 0.810 2.920 1.230 ;
        RECT  2.590 0.810 2.760 1.070 ;
        RECT  2.465 1.815 2.625 2.405 ;
        RECT  2.365 1.815 2.465 2.075 ;
        RECT  2.185 2.585 2.355 2.765 ;
        RECT  2.025 1.860 2.185 2.765 ;
        RECT  1.925 2.945 2.185 3.205 ;
        RECT  1.720 1.860 2.025 2.020 ;
        RECT  0.125 2.605 2.025 2.765 ;
        RECT  0.555 2.945 1.925 3.105 ;
        RECT  1.720 0.790 1.875 1.050 ;
        RECT  1.365 2.265 1.845 2.425 ;
        RECT  1.560 0.790 1.720 2.020 ;
        RECT  1.205 1.035 1.365 2.425 ;
        RECT  1.105 1.035 1.205 1.295 ;
        RECT  0.325 2.265 1.205 2.425 ;
        RECT  0.285 2.945 0.555 3.160 ;
        RECT  0.325 0.975 0.400 1.235 ;
        RECT  0.165 0.975 0.325 2.425 ;
        RECT  0.140 0.975 0.165 1.235 ;
    END
END EDFFHQX8

MACRO EDFFHQX4
    CLASS CORE ;
    FOREIGN EDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.560 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.925 0.695 15.975 2.585 ;
        RECT  15.665 0.600 15.925 3.070 ;
        END
        ANTENNADIFFAREA     0.7980 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 1.695 3.125 1.955 ;
        RECT  3.045 1.695 3.095 1.990 ;
        RECT  2.885 1.410 3.045 1.990 ;
        RECT  2.540 1.410 2.885 1.570 ;
        RECT  2.380 0.585 2.540 1.570 ;
        RECT  2.130 0.585 2.380 0.745 ;
        RECT  1.870 0.585 2.130 0.855 ;
        END
        ANTENNAGATEAREA     0.2626 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.150 0.920 1.985 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.160 6.300 1.420 ;
        RECT  5.645 1.160 5.855 1.580 ;
        RECT  5.360 1.160 5.645 1.420 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.435 -0.250 16.560 0.250 ;
        RECT  16.175 -0.250 16.435 1.115 ;
        RECT  15.385 -0.250 16.175 0.250 ;
        RECT  15.125 -0.250 15.385 0.405 ;
        RECT  14.535 -0.250 15.125 0.250 ;
        RECT  14.275 -0.250 14.535 0.405 ;
        RECT  5.455 -0.250 14.275 0.250 ;
        RECT  5.195 -0.250 5.455 0.405 ;
        RECT  4.330 -0.250 5.195 0.250 ;
        RECT  4.070 -0.250 4.330 0.405 ;
        RECT  2.350 -0.250 4.070 0.250 ;
        RECT  2.090 -0.250 2.350 0.405 ;
        RECT  0.810 -0.250 2.090 0.250 ;
        RECT  0.550 -0.250 0.810 0.405 ;
        RECT  0.000 -0.250 0.550 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.435 3.440 16.560 3.940 ;
        RECT  16.175 2.275 16.435 3.940 ;
        RECT  15.410 3.440 16.175 3.940 ;
        RECT  15.150 2.955 15.410 3.940 ;
        RECT  14.390 3.440 15.150 3.940 ;
        RECT  14.130 3.285 14.390 3.940 ;
        RECT  11.835 3.440 14.130 3.940 ;
        RECT  11.575 3.285 11.835 3.940 ;
        RECT  10.755 3.440 11.575 3.940 ;
        RECT  10.495 3.285 10.755 3.940 ;
        RECT  9.485 3.440 10.495 3.940 ;
        RECT  9.225 2.890 9.485 3.940 ;
        RECT  7.775 3.440 9.225 3.940 ;
        RECT  7.515 3.285 7.775 3.940 ;
        RECT  6.685 3.440 7.515 3.940 ;
        RECT  6.425 3.285 6.685 3.940 ;
        RECT  4.735 3.440 6.425 3.940 ;
        RECT  4.475 3.285 4.735 3.940 ;
        RECT  2.795 3.440 4.475 3.940 ;
        RECT  2.535 3.285 2.795 3.940 ;
        RECT  1.375 3.440 2.535 3.940 ;
        RECT  1.115 3.285 1.375 3.940 ;
        RECT  0.000 3.440 1.115 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.380 1.490 15.480 1.750 ;
        RECT  15.220 1.490 15.380 2.775 ;
        RECT  13.315 2.615 15.220 2.775 ;
        RECT  14.915 1.035 15.015 1.295 ;
        RECT  14.915 2.175 15.015 2.435 ;
        RECT  14.755 1.035 14.915 2.435 ;
        RECT  14.025 1.035 14.755 1.195 ;
        RECT  14.125 1.555 14.755 1.820 ;
        RECT  13.865 0.470 14.025 1.195 ;
        RECT  10.440 0.470 13.865 0.630 ;
        RECT  13.645 1.375 13.805 2.350 ;
        RECT  13.430 3.060 13.690 3.260 ;
        RECT  13.145 0.810 13.685 1.085 ;
        RECT  13.495 1.375 13.645 1.535 ;
        RECT  13.335 1.265 13.495 1.535 ;
        RECT  12.175 3.060 13.430 3.220 ;
        RECT  13.145 2.280 13.315 2.880 ;
        RECT  13.055 0.810 13.145 2.880 ;
        RECT  12.985 0.810 13.055 2.760 ;
        RECT  11.925 0.810 12.985 0.970 ;
        RECT  12.360 2.600 12.985 2.760 ;
        RECT  12.705 2.125 12.805 2.385 ;
        RECT  12.705 1.150 12.745 1.310 ;
        RECT  12.545 1.150 12.705 2.385 ;
        RECT  11.745 1.150 12.545 1.310 ;
        RECT  11.295 2.160 12.545 2.320 ;
        RECT  12.295 2.550 12.360 2.760 ;
        RECT  12.035 2.500 12.295 2.760 ;
        RECT  12.015 2.940 12.175 3.220 ;
        RECT  11.405 1.490 12.155 1.650 ;
        RECT  9.925 2.940 12.015 3.100 ;
        RECT  11.585 0.870 11.745 1.310 ;
        RECT  11.015 0.870 11.585 1.030 ;
        RECT  11.245 1.240 11.405 1.650 ;
        RECT  11.035 2.125 11.295 2.725 ;
        RECT  10.835 1.240 11.245 1.400 ;
        RECT  10.495 1.585 11.065 1.845 ;
        RECT  10.265 2.410 11.035 2.570 ;
        RECT  10.675 0.810 10.835 1.400 ;
        RECT  10.100 0.810 10.675 0.970 ;
        RECT  10.335 1.150 10.495 2.180 ;
        RECT  10.280 0.440 10.440 0.630 ;
        RECT  8.455 1.150 10.335 1.310 ;
        RECT  9.845 2.020 10.335 2.180 ;
        RECT  9.660 0.440 10.280 0.600 ;
        RECT  9.840 0.780 10.100 0.970 ;
        RECT  9.765 2.550 9.925 3.100 ;
        RECT  9.585 2.020 9.845 2.315 ;
        RECT  7.475 0.810 9.840 0.970 ;
        RECT  9.030 2.550 9.765 2.710 ;
        RECT  9.500 0.440 9.660 0.630 ;
        RECT  9.360 1.555 9.620 1.815 ;
        RECT  8.625 2.020 9.585 2.180 ;
        RECT  5.795 0.470 9.500 0.630 ;
        RECT  8.185 1.555 9.360 1.715 ;
        RECT  8.870 2.550 9.030 2.765 ;
        RECT  8.185 2.605 8.870 2.765 ;
        RECT  8.195 2.945 8.795 3.215 ;
        RECT  8.365 2.020 8.625 2.405 ;
        RECT  3.960 2.945 8.195 3.105 ;
        RECT  8.025 1.245 8.185 2.765 ;
        RECT  7.945 1.245 8.025 1.410 ;
        RECT  4.300 2.605 8.025 2.765 ;
        RECT  7.685 1.150 7.945 1.410 ;
        RECT  7.475 1.650 7.845 1.910 ;
        RECT  7.315 0.810 7.475 2.290 ;
        RECT  6.915 0.830 7.315 1.090 ;
        RECT  7.235 2.130 7.315 2.290 ;
        RECT  6.975 2.130 7.235 2.390 ;
        RECT  6.710 1.650 7.065 1.935 ;
        RECT  5.615 2.230 6.975 2.390 ;
        RECT  6.550 0.810 6.710 1.935 ;
        RECT  5.975 0.810 6.550 0.970 ;
        RECT  5.395 1.775 6.550 1.935 ;
        RECT  5.635 0.470 5.795 0.970 ;
        RECT  5.180 0.810 5.635 0.970 ;
        RECT  5.135 1.775 5.395 2.060 ;
        RECT  5.020 0.810 5.180 1.320 ;
        RECT  4.745 1.160 5.020 1.320 ;
        RECT  4.740 0.555 4.840 0.815 ;
        RECT  4.485 1.160 4.745 1.420 ;
        RECT  4.580 0.555 4.740 0.870 ;
        RECT  4.300 0.710 4.580 0.870 ;
        RECT  4.140 0.710 4.300 2.765 ;
        RECT  3.800 0.645 3.960 3.105 ;
        RECT  3.440 0.645 3.800 0.805 ;
        RECT  3.675 2.200 3.800 2.800 ;
        RECT  3.625 2.530 3.675 2.800 ;
        RECT  2.435 2.530 3.625 2.690 ;
        RECT  3.465 0.985 3.595 1.245 ;
        RECT  3.435 0.985 3.465 2.350 ;
        RECT  3.180 0.545 3.440 0.805 ;
        RECT  3.305 1.030 3.435 2.350 ;
        RECT  2.880 1.030 3.305 1.190 ;
        RECT  2.705 2.190 3.305 2.350 ;
        RECT  2.720 0.820 2.880 1.190 ;
        RECT  2.545 1.815 2.705 2.350 ;
        RECT  2.485 1.815 2.545 2.075 ;
        RECT  2.305 2.530 2.435 2.765 ;
        RECT  2.145 1.920 2.305 2.765 ;
        RECT  2.005 2.945 2.265 3.205 ;
        RECT  1.890 1.920 2.145 2.080 ;
        RECT  0.205 2.605 2.145 2.765 ;
        RECT  0.695 2.945 2.005 3.105 ;
        RECT  1.890 1.035 1.990 1.295 ;
        RECT  1.360 2.265 1.925 2.425 ;
        RECT  1.730 1.035 1.890 2.080 ;
        RECT  1.200 0.975 1.360 2.425 ;
        RECT  1.100 0.975 1.200 1.235 ;
        RECT  0.405 2.265 1.200 2.425 ;
        RECT  0.435 2.945 0.695 3.160 ;
        RECT  0.245 0.975 0.405 2.425 ;
        RECT  0.145 0.975 0.245 1.235 ;
    END
END EDFFHQX4

MACRO EDFFHQX2
    CLASS CORE ;
    FOREIGN EDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.875 0.600 10.915 2.585 ;
        RECT  10.655 0.600 10.875 3.050 ;
        RECT  10.615 1.955 10.655 3.050 ;
        END
        ANTENNADIFFAREA     0.7204 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 1.515 1.715 1.990 ;
        RECT  1.505 1.315 1.640 1.990 ;
        RECT  1.480 1.290 1.505 1.925 ;
        RECT  1.475 1.290 1.480 1.475 ;
        RECT  1.315 0.585 1.475 1.475 ;
        RECT  0.750 0.585 1.315 0.745 ;
        RECT  0.590 0.455 0.750 0.745 ;
        RECT  0.465 0.455 0.590 0.615 ;
        END
        ANTENNAGATEAREA     0.1495 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.535 1.400 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.410 4.175 1.995 ;
        RECT  3.785 1.640 4.015 1.995 ;
        END
        ANTENNAGATEAREA     0.2327 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.365 -0.250 11.040 0.250 ;
        RECT  9.425 -0.250 10.365 0.405 ;
        RECT  3.515 -0.250 9.425 0.250 ;
        RECT  3.255 -0.250 3.515 0.405 ;
        RECT  1.445 -0.250 3.255 0.250 ;
        RECT  1.185 -0.250 1.445 0.405 ;
        RECT  0.000 -0.250 1.185 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.315 3.440 11.040 3.940 ;
        RECT  10.055 3.285 10.315 3.940 ;
        RECT  9.495 3.440 10.055 3.940 ;
        RECT  9.235 2.890 9.495 3.940 ;
        RECT  7.110 3.440 9.235 3.940 ;
        RECT  6.850 3.285 7.110 3.940 ;
        RECT  5.710 3.440 6.850 3.940 ;
        RECT  5.450 3.285 5.710 3.940 ;
        RECT  3.675 3.440 5.450 3.940 ;
        RECT  3.415 3.285 3.675 3.940 ;
        RECT  1.785 3.440 3.415 3.940 ;
        RECT  1.625 3.075 1.785 3.940 ;
        RECT  0.000 3.440 1.625 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.275 1.050 10.435 2.285 ;
        RECT  9.480 1.050 10.275 1.210 ;
        RECT  9.885 2.125 10.275 2.285 ;
        RECT  9.105 1.625 10.095 1.785 ;
        RECT  9.625 2.125 9.885 2.385 ;
        RECT  9.445 2.125 9.625 2.315 ;
        RECT  9.320 0.585 9.480 1.210 ;
        RECT  9.285 2.055 9.445 2.315 ;
        RECT  8.630 0.585 9.320 0.745 ;
        RECT  8.945 0.925 9.105 2.655 ;
        RECT  8.380 0.925 8.945 1.085 ;
        RECT  8.550 2.495 8.945 2.655 ;
        RECT  8.550 2.945 8.810 3.245 ;
        RECT  8.605 2.055 8.765 2.315 ;
        RECT  8.470 0.470 8.630 0.745 ;
        RECT  8.385 1.265 8.605 1.525 ;
        RECT  8.385 2.055 8.605 2.215 ;
        RECT  8.290 2.495 8.550 2.755 ;
        RECT  6.780 2.945 8.550 3.105 ;
        RECT  7.080 0.470 8.470 0.630 ;
        RECT  8.225 1.265 8.385 2.215 ;
        RECT  8.200 1.265 8.225 1.425 ;
        RECT  8.040 0.810 8.200 1.425 ;
        RECT  6.735 0.810 8.040 0.970 ;
        RECT  7.880 1.605 8.040 2.750 ;
        RECT  7.860 1.605 7.880 1.765 ;
        RECT  7.780 2.150 7.880 2.750 ;
        RECT  7.700 1.150 7.860 1.765 ;
        RECT  7.010 2.420 7.780 2.580 ;
        RECT  7.595 1.150 7.700 1.310 ;
        RECT  7.415 1.645 7.520 1.940 ;
        RECT  7.255 1.300 7.415 2.240 ;
        RECT  6.535 1.300 7.255 1.460 ;
        RECT  6.440 2.080 7.255 2.240 ;
        RECT  6.920 0.430 7.080 0.630 ;
        RECT  6.295 0.430 6.920 0.590 ;
        RECT  6.620 2.605 6.780 3.105 ;
        RECT  6.475 0.780 6.735 0.970 ;
        RECT  6.095 1.640 6.735 1.900 ;
        RECT  6.095 2.605 6.620 2.765 ;
        RECT  6.325 1.150 6.535 1.460 ;
        RECT  5.275 0.810 6.475 0.970 ;
        RECT  6.280 2.080 6.440 2.340 ;
        RECT  6.275 1.150 6.325 1.310 ;
        RECT  6.135 0.430 6.295 0.630 ;
        RECT  6.235 3.100 6.285 3.260 ;
        RECT  6.025 2.945 6.235 3.260 ;
        RECT  4.015 0.470 6.135 0.630 ;
        RECT  5.935 1.270 6.095 2.765 ;
        RECT  2.815 2.945 6.025 3.105 ;
        RECT  5.615 1.270 5.935 1.430 ;
        RECT  3.355 2.605 5.935 2.765 ;
        RECT  5.275 1.650 5.755 1.910 ;
        RECT  5.455 1.170 5.615 1.430 ;
        RECT  5.115 0.810 5.275 2.385 ;
        RECT  4.735 0.810 5.115 0.970 ;
        RECT  4.215 2.225 5.115 2.385 ;
        RECT  4.515 1.650 4.935 1.940 ;
        RECT  4.355 0.870 4.515 2.040 ;
        RECT  4.225 0.870 4.355 1.030 ;
        RECT  3.855 0.470 4.015 0.760 ;
        RECT  3.825 0.600 3.855 0.760 ;
        RECT  3.665 0.600 3.825 1.425 ;
        RECT  3.345 1.265 3.665 1.425 ;
        RECT  3.325 0.820 3.485 1.080 ;
        RECT  3.195 1.715 3.355 2.765 ;
        RECT  3.185 1.265 3.345 1.525 ;
        RECT  3.005 0.920 3.325 1.080 ;
        RECT  3.005 1.715 3.195 1.875 ;
        RECT  2.845 0.920 3.005 1.875 ;
        RECT  2.815 2.375 2.915 2.635 ;
        RECT  2.665 2.055 2.815 3.105 ;
        RECT  2.655 0.920 2.665 3.105 ;
        RECT  2.505 0.920 2.655 2.215 ;
        RECT  1.445 2.735 2.655 2.895 ;
        RECT  2.425 0.920 2.505 1.080 ;
        RECT  2.265 0.435 2.425 1.080 ;
        RECT  2.275 2.395 2.405 2.555 ;
        RECT  2.275 1.260 2.325 1.520 ;
        RECT  2.115 1.260 2.275 2.555 ;
        RECT  1.985 0.435 2.265 0.595 ;
        RECT  2.055 1.260 2.115 1.420 ;
        RECT  1.105 2.395 2.115 2.555 ;
        RECT  1.895 0.945 2.055 1.420 ;
        RECT  1.655 0.945 1.895 1.105 ;
        RECT  1.285 2.735 1.445 3.220 ;
        RECT  1.135 2.005 1.290 2.165 ;
        RECT  0.385 3.060 1.285 3.220 ;
        RECT  0.975 0.945 1.135 2.165 ;
        RECT  0.945 2.395 1.105 2.875 ;
        RECT  0.635 0.945 0.975 1.105 ;
        RECT  0.285 0.895 0.385 1.155 ;
        RECT  0.285 2.360 0.385 3.220 ;
        RECT  0.225 0.895 0.285 3.220 ;
        RECT  0.125 0.895 0.225 2.960 ;
    END
END EDFFHQX2

MACRO EDFFHQX1
    CLASS CORE ;
    FOREIGN EDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.980 0.695 9.995 2.585 ;
        RECT  9.785 0.625 9.980 2.680 ;
        RECT  9.495 0.625 9.785 0.785 ;
        RECT  9.535 2.520 9.785 2.680 ;
        RECT  9.520 2.520 9.535 2.995 ;
        RECT  9.325 2.520 9.520 3.165 ;
        RECT  9.235 0.525 9.495 0.785 ;
        RECT  9.260 2.565 9.325 3.165 ;
        END
        ANTENNADIFFAREA     0.3638 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 0.470 1.795 0.905 ;
        END
        ANTENNAGATEAREA     0.1183 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.550 1.255 1.990 ;
        RECT  0.855 1.550 1.045 1.810 ;
        END
        ANTENNAGATEAREA     0.0923 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 1.290 3.625 1.690 ;
        END
        ANTENNAGATEAREA     0.1300 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.835 -0.250 10.120 0.250 ;
        RECT  8.575 -0.250 8.835 0.405 ;
        RECT  4.890 -0.250 8.575 0.250 ;
        RECT  4.290 -0.250 4.890 0.405 ;
        RECT  3.045 -0.250 4.290 0.250 ;
        RECT  2.785 -0.250 3.045 0.405 ;
        RECT  1.295 -0.250 2.785 0.250 ;
        RECT  1.035 -0.250 1.295 1.295 ;
        RECT  0.000 -0.250 1.035 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.955 3.440 10.120 3.940 ;
        RECT  8.695 2.615 8.955 3.940 ;
        RECT  7.020 3.440 8.695 3.940 ;
        RECT  6.760 3.285 7.020 3.940 ;
        RECT  4.845 3.440 6.760 3.940 ;
        RECT  4.585 3.285 4.845 3.940 ;
        RECT  3.180 3.440 4.585 3.940 ;
        RECT  2.920 3.285 3.180 3.940 ;
        RECT  1.455 3.440 2.920 3.940 ;
        RECT  1.195 3.115 1.455 3.940 ;
        RECT  0.000 3.440 1.195 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.490 1.035 9.590 1.295 ;
        RECT  9.490 2.025 9.550 2.335 ;
        RECT  9.330 1.035 9.490 2.335 ;
        RECT  9.040 1.035 9.330 1.195 ;
        RECT  9.290 2.025 9.330 2.335 ;
        RECT  8.700 2.175 9.290 2.335 ;
        RECT  8.990 1.405 9.150 1.665 ;
        RECT  8.880 0.720 9.040 1.195 ;
        RECT  8.700 1.405 8.990 1.565 ;
        RECT  8.330 0.720 8.880 0.880 ;
        RECT  8.540 1.065 8.700 1.565 ;
        RECT  8.540 1.885 8.700 2.335 ;
        RECT  8.020 1.065 8.540 1.225 ;
        RECT  8.200 1.405 8.360 3.100 ;
        RECT  8.170 0.470 8.330 0.880 ;
        RECT  7.590 2.940 8.200 3.100 ;
        RECT  5.230 0.470 8.170 0.630 ;
        RECT  7.990 1.065 8.020 2.005 ;
        RECT  7.925 0.965 7.990 2.005 ;
        RECT  7.860 0.965 7.925 2.725 ;
        RECT  7.830 0.965 7.860 1.225 ;
        RECT  7.765 1.845 7.860 2.725 ;
        RECT  7.720 2.120 7.765 2.725 ;
        RECT  7.650 1.405 7.680 1.665 ;
        RECT  7.490 0.810 7.650 1.665 ;
        RECT  7.330 2.940 7.590 3.215 ;
        RECT  5.570 0.810 7.490 0.970 ;
        RECT  7.310 2.135 7.420 2.760 ;
        RECT  5.875 2.940 7.330 3.100 ;
        RECT  7.150 1.150 7.310 2.760 ;
        RECT  6.390 2.600 7.150 2.760 ;
        RECT  6.810 1.635 6.970 1.930 ;
        RECT  6.485 1.635 6.810 1.895 ;
        RECT  6.325 1.180 6.485 2.420 ;
        RECT  5.750 1.180 6.325 1.340 ;
        RECT  5.565 2.260 6.325 2.420 ;
        RECT  5.385 1.815 6.145 2.075 ;
        RECT  5.715 2.605 5.875 3.100 ;
        RECT  5.385 2.605 5.715 2.765 ;
        RECT  5.410 0.810 5.570 1.085 ;
        RECT  5.275 2.945 5.535 3.260 ;
        RECT  4.890 0.925 5.410 1.085 ;
        RECT  5.225 1.265 5.385 2.765 ;
        RECT  4.390 2.945 5.275 3.105 ;
        RECT  5.070 0.470 5.230 0.745 ;
        RECT  5.070 1.265 5.225 1.425 ;
        RECT  4.045 2.605 5.225 2.765 ;
        RECT  2.720 0.585 5.070 0.745 ;
        RECT  4.970 1.730 5.045 1.990 ;
        RECT  4.890 1.730 4.970 2.405 ;
        RECT  4.810 0.925 4.890 2.405 ;
        RECT  4.730 0.925 4.810 1.890 ;
        RECT  3.615 2.245 4.810 2.405 ;
        RECT  4.390 0.925 4.730 1.085 ;
        RECT  4.140 1.450 4.550 1.710 ;
        RECT  4.230 2.945 4.390 3.260 ;
        RECT  3.600 3.100 4.230 3.260 ;
        RECT  3.980 0.950 4.140 2.035 ;
        RECT  3.785 2.605 4.045 2.920 ;
        RECT  3.880 0.950 3.980 1.110 ;
        RECT  3.660 1.875 3.980 2.035 ;
        RECT  3.060 2.605 3.785 2.765 ;
        RECT  3.060 0.950 3.630 1.110 ;
        RECT  3.440 2.945 3.600 3.260 ;
        RECT  2.390 2.945 3.440 3.105 ;
        RECT  2.900 0.950 3.060 2.765 ;
        RECT  2.560 0.585 2.720 1.720 ;
        RECT  2.365 2.150 2.390 3.105 ;
        RECT  2.230 0.625 2.365 3.105 ;
        RECT  2.205 0.625 2.230 2.930 ;
        RECT  2.175 0.625 2.205 0.785 ;
        RECT  1.015 2.770 2.205 2.930 ;
        RECT  1.975 0.525 2.175 0.785 ;
        RECT  1.835 1.610 2.025 1.870 ;
        RECT  1.835 1.085 1.935 1.245 ;
        RECT  1.820 2.050 1.925 2.310 ;
        RECT  1.820 1.085 1.835 1.870 ;
        RECT  1.660 1.085 1.820 2.590 ;
        RECT  0.675 2.430 1.660 2.590 ;
        RECT  0.855 2.770 1.015 3.125 ;
        RECT  0.335 2.965 0.855 3.125 ;
        RECT  0.675 1.990 0.845 2.250 ;
        RECT  0.675 1.035 0.785 1.295 ;
        RECT  0.515 1.035 0.675 2.250 ;
        RECT  0.515 2.430 0.675 2.785 ;
        RECT  0.335 0.455 0.385 0.715 ;
        RECT  0.175 0.455 0.335 3.125 ;
        RECT  0.125 0.455 0.175 0.715 ;
    END
END EDFFHQX1

MACRO DFFSRHQX8
    CLASS CORE ;
    FOREIGN DFFSRHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.560 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.290 4.800 1.745 ;
        END
        ANTENNAGATEAREA     0.2691 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.890 1.525 12.050 1.835 ;
        RECT  10.915 1.675 11.890 1.835 ;
        RECT  10.720 1.675 10.915 1.990 ;
        RECT  10.705 1.585 10.720 1.990 ;
        RECT  10.560 1.585 10.705 1.925 ;
        END
        ANTENNAGATEAREA     0.3419 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.910 1.105 15.975 2.585 ;
        RECT  15.650 0.595 15.910 3.045 ;
        RECT  15.305 0.935 15.650 2.435 ;
        RECT  14.890 0.935 15.305 1.275 ;
        RECT  14.890 2.105 15.305 2.435 ;
        RECT  14.630 0.595 14.890 1.275 ;
        RECT  14.630 2.105 14.890 3.045 ;
        END
        ANTENNADIFFAREA     1.6264 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.670 1.370 4.015 2.170 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.495 1.070 1.755 ;
        RECT  0.585 1.495 0.795 1.990 ;
        RECT  0.470 1.495 0.585 1.755 ;
        END
        ANTENNAGATEAREA     0.3783 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.420 -0.250 16.560 0.250 ;
        RECT  16.160 -0.250 16.420 1.095 ;
        RECT  15.400 -0.250 16.160 0.250 ;
        RECT  15.140 -0.250 15.400 0.755 ;
        RECT  14.350 -0.250 15.140 0.250 ;
        RECT  14.090 -0.250 14.350 0.405 ;
        RECT  12.635 -0.250 14.090 0.250 ;
        RECT  12.375 -0.250 12.635 0.405 ;
        RECT  9.890 -0.250 12.375 0.250 ;
        RECT  9.630 -0.250 9.890 0.405 ;
        RECT  7.645 -0.250 9.630 0.250 ;
        RECT  7.045 -0.250 7.645 0.405 ;
        RECT  5.215 -0.250 7.045 0.250 ;
        RECT  4.955 -0.250 5.215 0.405 ;
        RECT  3.515 -0.250 4.955 0.250 ;
        RECT  2.915 -0.250 3.515 0.405 ;
        RECT  1.270 -0.250 2.915 0.250 ;
        RECT  0.930 -0.250 1.270 0.405 ;
        RECT  0.670 -0.250 0.930 0.795 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.420 3.440 16.560 3.940 ;
        RECT  16.160 2.275 16.420 3.940 ;
        RECT  15.400 3.440 16.160 3.940 ;
        RECT  15.140 2.615 15.400 3.940 ;
        RECT  14.380 3.440 15.140 3.940 ;
        RECT  13.780 2.735 14.380 3.940 ;
        RECT  12.360 3.440 13.780 3.940 ;
        RECT  12.100 3.285 12.360 3.940 ;
        RECT  9.485 3.440 12.100 3.940 ;
        RECT  9.225 3.285 9.485 3.940 ;
        RECT  8.390 3.440 9.225 3.940 ;
        RECT  8.130 3.285 8.390 3.940 ;
        RECT  6.830 3.440 8.130 3.940 ;
        RECT  6.570 2.660 6.830 3.940 ;
        RECT  4.960 3.440 6.570 3.940 ;
        RECT  4.700 3.285 4.960 3.940 ;
        RECT  3.550 3.440 4.700 3.940 ;
        RECT  3.290 3.285 3.550 3.940 ;
        RECT  2.600 3.440 3.290 3.940 ;
        RECT  2.340 3.285 2.600 3.940 ;
        RECT  0.790 3.440 2.340 3.940 ;
        RECT  0.530 2.895 0.790 3.940 ;
        RECT  0.000 3.440 0.530 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.260 1.495 15.040 1.755 ;
        RECT  14.100 0.645 14.260 2.555 ;
        RECT  13.190 0.645 14.100 0.805 ;
        RECT  13.545 2.395 14.100 2.555 ;
        RECT  13.760 1.135 13.920 2.215 ;
        RECT  13.705 1.135 13.760 1.295 ;
        RECT  13.660 1.580 13.760 2.215 ;
        RECT  13.445 1.035 13.705 1.295 ;
        RECT  13.290 1.580 13.660 1.840 ;
        RECT  13.385 2.395 13.545 2.935 ;
        RECT  11.440 2.775 13.385 2.935 ;
        RECT  12.930 0.645 13.190 0.905 ;
        RECT  12.965 2.035 13.070 2.295 ;
        RECT  12.965 1.085 13.020 1.345 ;
        RECT  12.805 1.085 12.965 2.595 ;
        RECT  12.325 0.745 12.930 0.905 ;
        RECT  12.760 1.085 12.805 1.345 ;
        RECT  11.780 2.435 12.805 2.595 ;
        RECT  12.490 1.995 12.590 2.255 ;
        RECT  12.330 1.180 12.490 2.255 ;
        RECT  10.910 1.180 12.330 1.340 ;
        RECT  12.165 0.745 12.325 0.970 ;
        RECT  11.160 0.810 12.165 0.970 ;
        RECT  10.910 0.470 11.790 0.630 ;
        RECT  11.680 2.170 11.780 2.595 ;
        RECT  11.620 2.055 11.680 2.595 ;
        RECT  11.420 2.055 11.620 2.330 ;
        RECT  11.180 2.510 11.440 3.110 ;
        RECT  10.380 2.170 11.420 2.330 ;
        RECT  10.750 0.470 10.910 1.340 ;
        RECT  10.625 2.510 10.885 2.770 ;
        RECT  10.230 0.470 10.750 0.630 ;
        RECT  8.940 2.510 10.625 2.670 ;
        RECT  10.410 0.810 10.570 1.085 ;
        RECT  10.380 0.925 10.410 1.085 ;
        RECT  10.220 0.925 10.380 2.330 ;
        RECT  10.070 0.470 10.230 0.745 ;
        RECT  9.105 0.925 10.220 1.085 ;
        RECT  9.720 2.015 10.220 2.330 ;
        RECT  9.450 0.585 10.070 0.745 ;
        RECT  9.880 1.265 10.040 1.525 ;
        RECT  9.665 2.945 9.925 3.225 ;
        RECT  8.770 1.265 9.880 1.425 ;
        RECT  7.845 2.945 9.665 3.105 ;
        RECT  9.290 0.470 9.450 0.745 ;
        RECT  7.985 0.470 9.290 0.630 ;
        RECT  8.945 0.810 9.105 1.085 ;
        RECT  8.325 0.810 8.945 0.970 ;
        RECT  8.680 2.505 8.940 2.765 ;
        RECT  8.670 1.150 8.770 1.425 ;
        RECT  8.670 2.505 8.680 2.665 ;
        RECT  8.510 1.150 8.670 2.665 ;
        RECT  7.850 1.825 8.510 1.985 ;
        RECT  8.170 1.325 8.330 1.645 ;
        RECT  8.165 0.810 8.325 1.085 ;
        RECT  7.510 1.325 8.170 1.485 ;
        RECT  5.140 0.925 8.165 1.085 ;
        RECT  7.825 0.470 7.985 0.745 ;
        RECT  7.690 1.700 7.850 1.985 ;
        RECT  7.585 2.945 7.845 3.245 ;
        RECT  3.150 0.585 7.825 0.745 ;
        RECT  7.510 2.505 7.650 2.765 ;
        RECT  7.170 2.945 7.585 3.105 ;
        RECT  7.350 1.325 7.510 2.765 ;
        RECT  6.430 1.325 7.350 1.485 ;
        RECT  7.010 2.210 7.170 3.105 ;
        RECT  6.080 2.210 7.010 2.370 ;
        RECT  6.380 1.275 6.430 1.535 ;
        RECT  6.170 1.275 6.380 1.540 ;
        RECT  5.480 1.380 6.170 1.540 ;
        RECT  5.955 2.210 6.080 3.235 ;
        RECT  5.920 1.965 5.955 3.235 ;
        RECT  5.795 1.965 5.920 2.370 ;
        RECT  5.300 3.075 5.920 3.235 ;
        RECT  5.660 1.965 5.795 2.225 ;
        RECT  5.480 2.605 5.740 2.875 ;
        RECT  5.320 1.380 5.480 2.425 ;
        RECT  3.490 2.605 5.480 2.765 ;
        RECT  5.220 2.265 5.320 2.425 ;
        RECT  5.140 2.945 5.300 3.235 ;
        RECT  4.980 0.925 5.140 2.085 ;
        RECT  1.615 2.945 5.140 3.105 ;
        RECT  4.305 0.925 4.980 1.085 ;
        RECT  4.820 1.925 4.980 2.085 ;
        RECT  4.660 1.925 4.820 2.205 ;
        RECT  4.500 2.045 4.660 2.205 ;
        RECT  4.240 2.045 4.500 2.305 ;
        RECT  3.845 0.925 4.005 1.185 ;
        RECT  3.490 1.025 3.845 1.185 ;
        RECT  3.330 1.025 3.490 2.765 ;
        RECT  2.990 0.585 3.150 2.690 ;
        RECT  2.985 0.925 2.990 1.875 ;
        RECT  2.890 2.090 2.990 2.690 ;
        RECT  2.375 0.925 2.985 1.185 ;
        RECT  1.970 1.715 2.985 1.875 ;
        RECT  2.195 0.485 2.265 0.745 ;
        RECT  2.005 0.485 2.195 0.790 ;
        RECT  1.270 0.630 2.005 0.790 ;
        RECT  1.810 1.670 1.970 1.875 ;
        RECT  1.800 1.035 1.900 1.295 ;
        RECT  1.690 1.670 1.810 1.830 ;
        RECT  1.640 1.035 1.800 1.485 ;
        RECT  1.615 2.120 1.770 2.380 ;
        RECT  1.410 1.325 1.640 1.485 ;
        RECT  1.455 2.120 1.615 3.105 ;
        RECT  1.410 2.120 1.455 2.280 ;
        RECT  1.250 1.325 1.410 2.280 ;
        RECT  1.110 0.630 1.270 1.135 ;
        RECT  0.390 0.975 1.110 1.135 ;
        RECT  0.290 0.930 0.390 1.190 ;
        RECT  0.290 2.095 0.390 2.355 ;
        RECT  0.130 0.930 0.290 2.355 ;
    END
END DFFSRHQX8

MACRO DFFSRHQX4
    CLASS CORE ;
    FOREIGN DFFSRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.640 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.740 1.485 4.765 1.745 ;
        RECT  4.265 1.290 4.740 1.745 ;
        END
        ANTENNAGATEAREA     0.2691 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.840 1.520 12.100 1.835 ;
        RECT  10.915 1.675 11.840 1.835 ;
        RECT  10.720 1.675 10.915 1.990 ;
        RECT  10.705 1.535 10.720 1.990 ;
        RECT  10.560 1.535 10.705 1.835 ;
        END
        ANTENNAGATEAREA     0.3419 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.505 1.290 15.515 2.175 ;
        RECT  15.305 1.060 15.505 2.305 ;
        RECT  15.055 1.060 15.305 1.260 ;
        RECT  15.055 2.105 15.305 2.305 ;
        RECT  15.005 0.695 15.055 1.260 ;
        RECT  15.005 2.105 15.055 2.585 ;
        RECT  14.745 0.595 15.005 1.260 ;
        RECT  14.745 2.105 15.005 3.045 ;
        END
        ANTENNADIFFAREA     0.8132 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.670 1.370 4.015 2.170 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.495 1.070 1.755 ;
        RECT  0.585 1.495 0.795 1.990 ;
        RECT  0.470 1.495 0.585 1.755 ;
        END
        ANTENNAGATEAREA     0.3783 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.515 -0.250 15.640 0.250 ;
        RECT  15.255 -0.250 15.515 0.755 ;
        RECT  14.465 -0.250 15.255 0.250 ;
        RECT  13.865 -0.250 14.465 0.405 ;
        RECT  12.640 -0.250 13.865 0.250 ;
        RECT  12.380 -0.250 12.640 0.405 ;
        RECT  9.890 -0.250 12.380 0.250 ;
        RECT  9.630 -0.250 9.890 0.405 ;
        RECT  7.645 -0.250 9.630 0.250 ;
        RECT  7.045 -0.250 7.645 0.405 ;
        RECT  5.215 -0.250 7.045 0.250 ;
        RECT  4.955 -0.250 5.215 0.405 ;
        RECT  3.515 -0.250 4.955 0.250 ;
        RECT  2.915 -0.250 3.515 0.405 ;
        RECT  1.270 -0.250 2.915 0.250 ;
        RECT  0.930 -0.250 1.270 0.405 ;
        RECT  0.670 -0.250 0.930 0.795 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.515 3.440 15.640 3.940 ;
        RECT  15.255 2.615 15.515 3.940 ;
        RECT  14.495 3.440 15.255 3.940 ;
        RECT  13.895 2.955 14.495 3.940 ;
        RECT  12.360 3.440 13.895 3.940 ;
        RECT  12.100 3.285 12.360 3.940 ;
        RECT  9.485 3.440 12.100 3.940 ;
        RECT  9.225 3.285 9.485 3.940 ;
        RECT  8.390 3.440 9.225 3.940 ;
        RECT  8.130 3.285 8.390 3.940 ;
        RECT  6.830 3.440 8.130 3.940 ;
        RECT  6.570 2.660 6.830 3.940 ;
        RECT  4.960 3.440 6.570 3.940 ;
        RECT  4.700 3.285 4.960 3.940 ;
        RECT  3.550 3.440 4.700 3.940 ;
        RECT  3.290 3.285 3.550 3.940 ;
        RECT  2.600 3.440 3.290 3.940 ;
        RECT  2.340 3.285 2.600 3.940 ;
        RECT  0.790 3.440 2.340 3.940 ;
        RECT  0.530 2.895 0.790 3.940 ;
        RECT  0.000 3.440 0.530 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.330 1.495 15.040 1.755 ;
        RECT  14.170 0.695 14.330 2.580 ;
        RECT  13.190 0.695 14.170 0.855 ;
        RECT  14.100 1.495 14.170 1.755 ;
        RECT  13.545 2.420 14.170 2.580 ;
        RECT  13.760 1.135 13.920 2.215 ;
        RECT  13.705 1.135 13.760 1.295 ;
        RECT  13.660 1.580 13.760 2.215 ;
        RECT  13.445 1.035 13.705 1.295 ;
        RECT  13.245 1.580 13.660 1.840 ;
        RECT  13.385 2.420 13.545 2.935 ;
        RECT  11.440 2.775 13.385 2.935 ;
        RECT  12.930 0.645 13.190 0.905 ;
        RECT  12.875 1.085 13.020 1.345 ;
        RECT  12.875 2.035 13.020 2.295 ;
        RECT  12.535 0.745 12.930 0.905 ;
        RECT  12.715 1.085 12.875 2.595 ;
        RECT  11.825 2.435 12.715 2.595 ;
        RECT  12.375 0.745 12.535 1.000 ;
        RECT  12.375 1.180 12.535 2.210 ;
        RECT  11.160 0.840 12.375 1.000 ;
        RECT  10.910 1.180 12.375 1.340 ;
        RECT  12.275 2.050 12.375 2.210 ;
        RECT  11.680 2.170 11.825 2.595 ;
        RECT  10.910 0.470 11.795 0.630 ;
        RECT  11.665 2.055 11.680 2.595 ;
        RECT  11.420 2.055 11.665 2.330 ;
        RECT  11.180 2.510 11.440 3.110 ;
        RECT  10.380 2.170 11.420 2.330 ;
        RECT  10.750 0.470 10.910 1.340 ;
        RECT  10.625 2.605 10.885 2.865 ;
        RECT  10.230 0.470 10.750 0.630 ;
        RECT  8.940 2.605 10.625 2.765 ;
        RECT  10.410 0.810 10.570 1.085 ;
        RECT  10.380 0.925 10.410 1.085 ;
        RECT  10.220 0.925 10.380 2.330 ;
        RECT  10.070 0.470 10.230 0.745 ;
        RECT  9.105 0.925 10.220 1.085 ;
        RECT  9.975 2.070 10.220 2.330 ;
        RECT  9.450 0.585 10.070 0.745 ;
        RECT  9.880 1.265 10.040 1.530 ;
        RECT  9.665 2.945 9.925 3.260 ;
        RECT  8.770 1.370 9.880 1.530 ;
        RECT  7.845 2.945 9.665 3.105 ;
        RECT  9.290 0.470 9.450 0.745 ;
        RECT  7.985 0.470 9.290 0.630 ;
        RECT  8.945 0.810 9.105 1.085 ;
        RECT  8.325 0.810 8.945 0.970 ;
        RECT  8.680 2.505 8.940 2.765 ;
        RECT  8.670 1.150 8.770 1.530 ;
        RECT  8.670 2.505 8.680 2.665 ;
        RECT  8.510 1.150 8.670 2.665 ;
        RECT  7.850 1.825 8.510 1.985 ;
        RECT  8.170 1.325 8.330 1.645 ;
        RECT  8.165 0.810 8.325 1.085 ;
        RECT  7.510 1.325 8.170 1.485 ;
        RECT  5.110 0.925 8.165 1.085 ;
        RECT  7.825 0.470 7.985 0.745 ;
        RECT  7.690 1.700 7.850 1.985 ;
        RECT  7.585 2.945 7.845 3.245 ;
        RECT  3.150 0.585 7.825 0.745 ;
        RECT  7.510 2.505 7.650 2.765 ;
        RECT  7.170 2.945 7.585 3.105 ;
        RECT  7.350 1.325 7.510 2.765 ;
        RECT  6.430 1.325 7.350 1.485 ;
        RECT  7.010 2.210 7.170 3.105 ;
        RECT  6.080 2.210 7.010 2.370 ;
        RECT  6.380 1.275 6.430 1.535 ;
        RECT  6.170 1.275 6.380 1.540 ;
        RECT  5.480 1.380 6.170 1.540 ;
        RECT  5.955 2.210 6.080 3.235 ;
        RECT  5.920 1.965 5.955 3.235 ;
        RECT  5.795 1.965 5.920 2.370 ;
        RECT  5.300 3.075 5.920 3.235 ;
        RECT  5.660 1.965 5.795 2.225 ;
        RECT  5.480 2.605 5.740 2.875 ;
        RECT  5.320 1.380 5.480 2.425 ;
        RECT  3.490 2.605 5.480 2.765 ;
        RECT  5.220 2.265 5.320 2.425 ;
        RECT  5.140 2.945 5.300 3.235 ;
        RECT  1.615 2.945 5.140 3.105 ;
        RECT  5.005 0.925 5.110 2.085 ;
        RECT  4.950 0.925 5.005 2.205 ;
        RECT  4.305 0.925 4.950 1.085 ;
        RECT  4.845 1.925 4.950 2.205 ;
        RECT  4.500 2.045 4.845 2.205 ;
        RECT  4.240 2.045 4.500 2.305 ;
        RECT  3.845 0.925 4.005 1.185 ;
        RECT  3.490 1.025 3.845 1.185 ;
        RECT  3.330 1.025 3.490 2.765 ;
        RECT  2.990 0.585 3.150 2.690 ;
        RECT  2.985 0.925 2.990 1.875 ;
        RECT  2.890 2.090 2.990 2.690 ;
        RECT  2.375 0.925 2.985 1.185 ;
        RECT  2.055 1.715 2.985 1.875 ;
        RECT  2.195 0.485 2.265 0.745 ;
        RECT  2.005 0.485 2.195 0.790 ;
        RECT  1.795 1.620 2.055 1.880 ;
        RECT  1.275 0.630 2.005 0.790 ;
        RECT  1.640 1.035 1.900 1.295 ;
        RECT  1.615 2.120 1.770 2.380 ;
        RECT  1.615 1.135 1.640 1.295 ;
        RECT  1.455 1.135 1.615 3.105 ;
        RECT  1.115 0.630 1.275 1.190 ;
        RECT  0.390 1.030 1.115 1.190 ;
        RECT  0.290 0.930 0.390 1.190 ;
        RECT  0.290 2.095 0.390 2.355 ;
        RECT  0.130 0.930 0.290 2.355 ;
    END
END DFFSRHQX4

MACRO DFFSRHQX2
    CLASS CORE ;
    FOREIGN DFFSRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.340 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.615 1.290 4.015 1.840 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.645 1.825 9.905 2.085 ;
        RECT  9.535 1.825 9.645 1.990 ;
        RECT  9.325 1.700 9.535 1.990 ;
        RECT  8.285 1.830 9.325 1.990 ;
        END
        ANTENNAGATEAREA     0.2210 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.165 0.595 13.215 1.765 ;
        RECT  13.005 0.595 13.165 2.115 ;
        RECT  12.955 0.595 13.005 1.195 ;
        RECT  12.815 1.955 13.005 2.115 ;
        RECT  12.555 1.955 12.815 2.555 ;
        END
        ANTENNADIFFAREA     0.5653 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.665 1.290 3.095 1.845 ;
        RECT  2.615 1.295 2.665 1.455 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.835 1.920 ;
        RECT  0.575 1.660 0.585 1.920 ;
        END
        ANTENNAGATEAREA     0.2314 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.665 -0.250 13.340 0.250 ;
        RECT  12.405 -0.250 12.665 1.135 ;
        RECT  10.730 -0.250 12.405 0.250 ;
        RECT  10.470 -0.250 10.730 0.405 ;
        RECT  6.515 -0.250 10.470 0.250 ;
        RECT  6.255 -0.250 6.515 0.405 ;
        RECT  3.165 -0.250 6.255 0.250 ;
        RECT  2.225 -0.250 3.165 0.405 ;
        RECT  0.935 -0.250 2.225 0.250 ;
        RECT  0.675 -0.250 0.935 0.405 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.215 3.440 13.340 3.940 ;
        RECT  12.195 3.285 13.215 3.940 ;
        RECT  11.595 2.895 12.195 3.940 ;
        RECT  10.285 3.440 11.595 3.940 ;
        RECT  10.025 3.285 10.285 3.940 ;
        RECT  7.790 3.440 10.025 3.940 ;
        RECT  7.530 3.285 7.790 3.940 ;
        RECT  6.840 3.440 7.530 3.940 ;
        RECT  6.580 3.285 6.840 3.940 ;
        RECT  5.745 3.440 6.580 3.940 ;
        RECT  5.485 3.285 5.745 3.940 ;
        RECT  3.815 3.440 5.485 3.940 ;
        RECT  3.555 3.285 3.815 3.940 ;
        RECT  2.770 3.440 3.555 3.940 ;
        RECT  2.510 3.285 2.770 3.940 ;
        RECT  0.815 3.440 2.510 3.940 ;
        RECT  0.555 2.850 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.175 1.495 12.730 1.755 ;
        RECT  12.015 0.675 12.175 2.560 ;
        RECT  11.315 0.675 12.015 0.835 ;
        RECT  11.405 2.400 12.015 2.560 ;
        RECT  11.735 1.035 11.835 1.295 ;
        RECT  11.735 1.955 11.835 2.215 ;
        RECT  11.575 1.035 11.735 2.215 ;
        RECT  11.205 1.735 11.575 1.995 ;
        RECT  11.245 2.400 11.405 2.935 ;
        RECT  11.215 0.625 11.315 0.885 ;
        RECT  9.335 2.775 11.245 2.935 ;
        RECT  11.055 0.625 11.215 1.080 ;
        RECT  10.950 1.300 11.115 1.460 ;
        RECT  9.505 0.920 11.055 1.080 ;
        RECT  10.950 2.045 10.985 2.305 ;
        RECT  10.885 1.300 10.950 2.305 ;
        RECT  10.790 1.300 10.885 2.595 ;
        RECT  10.725 2.045 10.790 2.595 ;
        RECT  9.595 2.435 10.725 2.595 ;
        RECT  10.285 2.095 10.505 2.255 ;
        RECT  10.125 1.360 10.285 2.255 ;
        RECT  9.065 1.360 10.125 1.520 ;
        RECT  9.335 2.265 9.595 2.595 ;
        RECT  9.245 0.920 9.505 1.180 ;
        RECT  9.065 0.470 9.455 0.630 ;
        RECT  8.085 2.265 9.335 2.425 ;
        RECT  9.075 2.775 9.335 3.105 ;
        RECT  8.905 0.470 9.065 1.520 ;
        RECT  6.860 0.470 8.905 0.630 ;
        RECT  8.565 2.605 8.825 2.895 ;
        RECT  8.550 0.810 8.710 1.650 ;
        RECT  7.390 2.605 8.565 2.765 ;
        RECT  8.130 3.100 8.565 3.260 ;
        RECT  7.200 0.810 8.550 0.970 ;
        RECT  8.085 1.490 8.550 1.650 ;
        RECT  7.540 1.150 8.370 1.310 ;
        RECT  7.970 2.945 8.130 3.260 ;
        RECT  7.925 1.490 8.085 2.425 ;
        RECT  6.300 2.945 7.970 3.105 ;
        RECT  7.805 2.020 7.925 2.280 ;
        RECT  7.380 1.150 7.540 1.425 ;
        RECT  7.230 2.135 7.390 2.765 ;
        RECT  6.965 1.265 7.380 1.425 ;
        RECT  7.130 2.135 7.230 2.395 ;
        RECT  7.040 0.810 7.200 1.085 ;
        RECT  6.965 2.135 7.130 2.295 ;
        RECT  5.735 0.925 7.040 1.085 ;
        RECT  6.805 1.265 6.965 2.295 ;
        RECT  6.700 0.470 6.860 0.745 ;
        RECT  6.515 1.265 6.805 1.425 ;
        RECT  6.355 1.935 6.805 2.195 ;
        RECT  6.075 0.585 6.700 0.745 ;
        RECT  6.175 1.455 6.335 1.715 ;
        RECT  6.040 2.925 6.300 3.185 ;
        RECT  5.395 1.505 6.175 1.665 ;
        RECT  5.845 2.485 6.105 2.745 ;
        RECT  5.915 0.470 6.075 0.745 ;
        RECT  5.950 2.925 6.040 3.105 ;
        RECT  5.055 2.925 5.950 3.085 ;
        RECT  3.505 0.470 5.915 0.630 ;
        RECT  5.395 2.485 5.845 2.645 ;
        RECT  5.575 0.810 5.735 1.085 ;
        RECT  3.845 0.810 5.575 0.970 ;
        RECT  5.235 1.150 5.395 2.645 ;
        RECT  4.355 1.150 5.235 1.310 ;
        RECT  4.965 1.655 5.055 3.085 ;
        RECT  4.895 1.655 4.965 3.260 ;
        RECT  4.695 1.655 4.895 1.815 ;
        RECT  4.805 2.925 4.895 3.260 ;
        RECT  4.185 3.100 4.805 3.260 ;
        RECT  4.455 2.090 4.715 2.350 ;
        RECT  4.535 1.555 4.695 1.815 ;
        RECT  4.365 2.605 4.625 2.910 ;
        RECT  4.355 2.090 4.455 2.250 ;
        RECT  3.205 2.605 4.365 2.765 ;
        RECT  4.195 1.150 4.355 2.250 ;
        RECT  4.025 2.945 4.185 3.260 ;
        RECT  1.795 2.945 4.025 3.105 ;
        RECT  3.685 0.810 3.845 1.110 ;
        RECT  3.435 0.950 3.685 1.110 ;
        RECT  3.345 0.470 3.505 0.745 ;
        RECT  3.275 0.950 3.435 2.185 ;
        RECT  1.970 0.585 3.345 0.745 ;
        RECT  3.170 0.950 3.275 1.110 ;
        RECT  3.235 2.025 3.275 2.185 ;
        RECT  2.975 2.025 3.235 2.285 ;
        RECT  2.945 2.585 3.205 2.765 ;
        RECT  2.485 2.605 2.945 2.765 ;
        RECT  2.310 0.925 2.920 1.085 ;
        RECT  2.325 1.620 2.485 2.765 ;
        RECT  2.310 1.620 2.325 1.780 ;
        RECT  2.150 0.925 2.310 1.780 ;
        RECT  1.970 1.960 2.145 2.220 ;
        RECT  1.810 0.585 1.970 2.220 ;
        RECT  1.675 0.815 1.810 1.075 ;
        RECT  1.365 1.870 1.810 2.130 ;
        RECT  1.635 2.615 1.795 3.105 ;
        RECT  1.535 2.615 1.635 2.875 ;
        RECT  1.175 2.615 1.535 2.775 ;
        RECT  1.235 0.620 1.495 0.880 ;
        RECT  1.175 1.065 1.365 1.225 ;
        RECT  0.385 0.720 1.235 0.880 ;
        RECT  1.015 1.065 1.175 2.775 ;
        RECT  0.225 0.720 0.385 2.365 ;
        RECT  0.125 1.030 0.225 1.290 ;
        RECT  0.125 2.105 0.225 2.365 ;
    END
END DFFSRHQX2

MACRO DFFSRHQX1
    CLASS CORE ;
    FOREIGN DFFSRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.420 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.290 3.210 1.940 ;
        END
        ANTENNAGATEAREA     0.1365 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.075 1.755 9.665 1.915 ;
        RECT  8.435 1.615 9.075 1.990 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.245 1.105 12.295 2.615 ;
        RECT  12.110 0.915 12.245 2.615 ;
        RECT  12.085 0.815 12.110 2.615 ;
        RECT  11.840 0.815 12.085 1.075 ;
        RECT  12.035 2.015 12.085 2.615 ;
        END
        ANTENNADIFFAREA     0.3944 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.345 1.290 2.635 1.940 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 1.290 0.795 1.845 ;
        RECT  0.530 1.585 0.545 1.845 ;
        END
        ANTENNAGATEAREA     0.1456 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.550 -0.250 12.420 0.250 ;
        RECT  11.290 -0.250 11.550 0.405 ;
        RECT  10.100 -0.250 11.290 0.250 ;
        RECT  9.840 -0.250 10.100 0.405 ;
        RECT  7.080 -0.250 9.840 0.250 ;
        RECT  6.140 -0.250 7.080 0.405 ;
        RECT  3.835 -0.250 6.140 0.250 ;
        RECT  3.575 -0.250 3.835 0.405 ;
        RECT  2.385 -0.250 3.575 0.250 ;
        RECT  2.125 -0.250 2.385 0.405 ;
        RECT  0.965 -0.250 2.125 0.250 ;
        RECT  0.705 -0.250 0.965 0.405 ;
        RECT  0.000 -0.250 0.705 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.745 3.440 12.420 3.940 ;
        RECT  11.485 2.780 11.745 3.940 ;
        RECT  9.970 3.440 11.485 3.940 ;
        RECT  9.710 3.285 9.970 3.940 ;
        RECT  7.615 3.440 9.710 3.940 ;
        RECT  7.355 3.285 7.615 3.940 ;
        RECT  6.585 3.440 7.355 3.940 ;
        RECT  5.645 3.285 6.585 3.940 ;
        RECT  4.035 3.440 5.645 3.940 ;
        RECT  3.775 3.285 4.035 3.940 ;
        RECT  2.515 3.440 3.775 3.940 ;
        RECT  2.255 3.285 2.515 3.940 ;
        RECT  0.795 3.440 2.255 3.940 ;
        RECT  0.535 2.555 0.795 3.940 ;
        RECT  0.000 3.440 0.535 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.590 1.255 11.690 2.595 ;
        RECT  11.530 0.585 11.590 2.595 ;
        RECT  11.430 0.585 11.530 1.515 ;
        RECT  9.860 2.435 11.530 2.595 ;
        RECT  10.680 0.585 11.430 0.745 ;
        RECT  11.070 1.960 11.320 2.220 ;
        RECT  10.910 0.955 11.070 2.220 ;
        RECT  10.420 0.430 10.680 0.745 ;
        RECT  10.540 1.705 10.640 1.965 ;
        RECT  10.380 0.930 10.540 2.255 ;
        RECT  8.935 0.585 10.420 0.745 ;
        RECT  10.255 0.930 10.380 1.090 ;
        RECT  9.415 2.095 10.380 2.255 ;
        RECT  10.060 1.755 10.160 1.915 ;
        RECT  9.900 1.275 10.060 1.915 ;
        RECT  8.595 1.275 9.900 1.435 ;
        RECT  9.700 2.435 9.860 3.075 ;
        RECT  8.815 2.915 9.700 3.075 ;
        RECT  9.255 2.095 9.415 2.565 ;
        RECT  9.020 2.265 9.255 2.565 ;
        RECT  8.255 2.265 9.020 2.425 ;
        RECT  8.775 0.585 8.935 1.095 ;
        RECT  8.435 0.585 8.595 1.435 ;
        RECT  5.400 0.585 8.435 0.745 ;
        RECT  8.175 2.605 8.435 2.865 ;
        RECT  8.095 0.925 8.255 2.425 ;
        RECT  7.955 3.100 8.250 3.260 ;
        RECT  7.315 2.605 8.175 2.765 ;
        RECT  3.550 0.925 8.095 1.085 ;
        RECT  7.755 2.265 8.095 2.425 ;
        RECT  7.795 2.945 7.955 3.260 ;
        RECT  7.315 1.265 7.915 1.425 ;
        RECT  5.055 2.945 7.795 3.105 ;
        RECT  7.495 2.095 7.755 2.425 ;
        RECT  7.155 1.265 7.315 2.765 ;
        RECT  6.175 1.265 7.155 1.425 ;
        RECT  6.495 2.605 7.155 2.765 ;
        RECT  6.855 2.165 6.975 2.425 ;
        RECT  6.695 1.760 6.855 2.425 ;
        RECT  6.055 1.760 6.695 1.920 ;
        RECT  6.335 2.185 6.495 2.765 ;
        RECT  6.235 2.185 6.335 2.445 ;
        RECT  5.895 1.760 6.055 2.765 ;
        RECT  5.495 1.760 5.895 1.920 ;
        RECT  5.555 2.605 5.895 2.765 ;
        RECT  5.055 2.165 5.715 2.425 ;
        RECT  5.335 1.265 5.495 1.920 ;
        RECT  5.140 0.560 5.400 0.745 ;
        RECT  3.890 1.265 5.335 1.425 ;
        RECT  1.825 0.585 5.140 0.745 ;
        RECT  4.895 1.695 5.055 3.245 ;
        RECT  4.140 1.695 4.895 1.855 ;
        RECT  4.375 3.085 4.895 3.245 ;
        RECT  4.555 2.605 4.715 2.905 ;
        RECT  3.890 2.265 4.595 2.425 ;
        RECT  3.255 2.605 4.555 2.765 ;
        RECT  4.215 2.945 4.375 3.245 ;
        RECT  3.595 2.945 4.215 3.105 ;
        RECT  3.730 1.265 3.890 2.425 ;
        RECT  3.435 2.945 3.595 3.245 ;
        RECT  3.390 0.925 3.550 2.345 ;
        RECT  2.865 3.085 3.435 3.245 ;
        RECT  3.145 0.925 3.390 1.110 ;
        RECT  3.025 2.185 3.390 2.345 ;
        RECT  3.095 2.605 3.255 2.905 ;
        RECT  2.845 2.605 3.095 2.765 ;
        RECT  2.165 0.925 2.895 1.085 ;
        RECT  2.705 2.945 2.865 3.245 ;
        RECT  2.685 2.130 2.845 2.765 ;
        RECT  1.685 2.945 2.705 3.105 ;
        RECT  2.165 2.130 2.685 2.290 ;
        RECT  1.935 2.470 2.195 2.730 ;
        RECT  2.005 0.925 2.165 2.290 ;
        RECT  1.825 2.470 1.935 2.630 ;
        RECT  1.665 0.445 1.825 2.630 ;
        RECT  1.425 2.810 1.685 3.105 ;
        RECT  1.415 1.650 1.665 1.920 ;
        RECT  1.295 0.645 1.455 0.905 ;
        RECT  1.235 2.810 1.425 2.970 ;
        RECT  1.235 1.085 1.395 1.245 ;
        RECT  0.385 0.745 1.295 0.905 ;
        RECT  1.075 1.085 1.235 2.970 ;
        RECT  0.335 0.745 0.385 1.110 ;
        RECT  0.335 2.030 0.385 2.290 ;
        RECT  0.175 0.745 0.335 2.290 ;
        RECT  0.125 0.850 0.175 1.110 ;
        RECT  0.125 2.030 0.175 2.290 ;
    END
END DFFSRHQX1

MACRO DFFSHQX8
    CLASS CORE ;
    FOREIGN DFFSHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.560 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.660 1.700 8.155 2.085 ;
        END
        ANTENNAGATEAREA     0.3510 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.860 1.515 15.975 1.765 ;
        RECT  15.600 0.595 15.860 3.060 ;
        RECT  14.840 1.700 15.600 2.400 ;
        RECT  14.580 0.775 14.840 3.060 ;
        END
        ANTENNADIFFAREA     1.6234 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.620 3.715 1.990 ;
        RECT  3.210 1.700 3.220 1.980 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.495 1.930 1.755 ;
        RECT  1.485 1.495 1.715 1.990 ;
        RECT  0.990 1.495 1.485 1.755 ;
        END
        ANTENNAGATEAREA     0.4563 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.370 -0.250 16.560 0.250 ;
        RECT  16.110 -0.250 16.370 1.095 ;
        RECT  15.350 -0.250 16.110 0.250 ;
        RECT  15.090 -0.250 15.350 1.095 ;
        RECT  14.440 -0.250 15.090 0.250 ;
        RECT  14.180 -0.250 14.440 0.405 ;
        RECT  12.300 -0.250 14.180 0.250 ;
        RECT  12.660 1.000 12.920 1.260 ;
        RECT  12.300 1.000 12.660 1.160 ;
        RECT  12.140 -0.250 12.300 1.160 ;
        RECT  9.980 -0.250 12.140 0.250 ;
        RECT  9.720 -0.250 9.980 0.575 ;
        RECT  8.895 -0.250 9.720 0.250 ;
        RECT  8.635 -0.250 8.895 0.575 ;
        RECT  8.325 -0.250 8.635 0.250 ;
        RECT  8.065 -0.250 8.325 0.575 ;
        RECT  7.225 -0.250 8.065 0.250 ;
        RECT  6.965 -0.250 7.225 0.625 ;
        RECT  4.030 -0.250 6.965 0.250 ;
        RECT  3.770 -0.250 4.030 0.405 ;
        RECT  2.535 -0.250 3.770 0.250 ;
        RECT  2.275 -0.250 2.535 1.065 ;
        RECT  1.020 -0.250 2.275 0.250 ;
        RECT  0.760 -0.250 1.020 0.405 ;
        RECT  0.000 -0.250 0.760 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.370 3.440 16.560 3.940 ;
        RECT  16.110 2.275 16.370 3.940 ;
        RECT  15.350 3.440 16.110 3.940 ;
        RECT  15.090 2.615 15.350 3.940 ;
        RECT  14.090 3.440 15.090 3.940 ;
        RECT  13.830 3.285 14.090 3.940 ;
        RECT  11.890 3.440 13.830 3.940 ;
        RECT  11.630 3.285 11.890 3.940 ;
        RECT  9.285 3.440 11.630 3.940 ;
        RECT  9.025 2.955 9.285 3.940 ;
        RECT  7.675 3.440 9.025 3.940 ;
        RECT  7.415 3.285 7.675 3.940 ;
        RECT  6.605 3.440 7.415 3.940 ;
        RECT  6.345 3.285 6.605 3.940 ;
        RECT  4.620 3.440 6.345 3.940 ;
        RECT  4.360 3.285 4.620 3.940 ;
        RECT  3.530 3.440 4.360 3.940 ;
        RECT  3.270 3.285 3.530 3.940 ;
        RECT  1.670 3.440 3.270 3.940 ;
        RECT  1.410 3.285 1.670 3.940 ;
        RECT  0.000 3.440 1.410 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.210 0.590 14.370 3.105 ;
        RECT  14.000 0.590 14.210 0.750 ;
        RECT  13.420 2.945 14.210 3.105 ;
        RECT  13.930 1.640 14.030 2.750 ;
        RECT  13.840 0.470 14.000 0.750 ;
        RECT  13.870 0.930 13.930 2.750 ;
        RECT  13.770 0.930 13.870 1.900 ;
        RECT  13.080 2.590 13.870 2.750 ;
        RECT  12.660 0.470 13.840 0.630 ;
        RECT  13.660 0.930 13.770 1.090 ;
        RECT  13.390 2.250 13.690 2.410 ;
        RECT  13.500 0.810 13.660 1.090 ;
        RECT  13.400 0.810 13.500 0.970 ;
        RECT  13.390 1.270 13.490 1.530 ;
        RECT  13.260 2.945 13.420 3.260 ;
        RECT  13.230 1.270 13.390 2.410 ;
        RECT  12.790 3.100 13.260 3.260 ;
        RECT  12.305 1.765 13.230 1.925 ;
        RECT  12.920 2.590 13.080 2.865 ;
        RECT  11.625 2.705 12.920 2.865 ;
        RECT  12.480 2.265 12.740 2.525 ;
        RECT  11.965 2.265 12.480 2.425 ;
        RECT  12.145 1.765 12.305 2.045 ;
        RECT  11.900 1.555 11.965 2.425 ;
        RECT  11.805 0.470 11.900 2.425 ;
        RECT  11.740 0.470 11.805 1.715 ;
        RECT  10.320 0.470 11.740 0.630 ;
        RECT  11.560 1.905 11.625 2.865 ;
        RECT  11.465 0.810 11.560 2.865 ;
        RECT  11.400 0.810 11.465 2.065 ;
        RECT  10.660 0.810 11.400 0.970 ;
        RECT  10.825 1.905 11.400 2.065 ;
        RECT  11.125 2.275 11.285 3.220 ;
        RECT  10.345 3.060 11.125 3.220 ;
        RECT  11.000 1.155 11.100 1.315 ;
        RECT  10.840 1.155 11.000 1.725 ;
        RECT  10.345 1.565 10.840 1.725 ;
        RECT  10.665 1.905 10.825 2.880 ;
        RECT  10.565 2.280 10.665 2.880 ;
        RECT  10.500 0.810 10.660 1.315 ;
        RECT  10.205 1.155 10.500 1.315 ;
        RECT  10.185 1.565 10.345 3.220 ;
        RECT  10.205 0.470 10.320 0.915 ;
        RECT  10.160 0.470 10.205 0.945 ;
        RECT  9.860 2.165 10.185 2.425 ;
        RECT  9.945 0.755 10.160 0.945 ;
        RECT  9.845 2.615 10.005 3.215 ;
        RECT  7.785 0.755 9.945 0.915 ;
        RECT  9.755 1.250 9.860 2.425 ;
        RECT  8.565 2.615 9.845 2.775 ;
        RECT  9.700 1.095 9.755 2.425 ;
        RECT  9.595 1.095 9.700 1.410 ;
        RECT  9.535 2.165 9.700 2.425 ;
        RECT  9.175 1.095 9.595 1.255 ;
        RECT  8.775 2.265 9.535 2.425 ;
        RECT  8.920 1.590 9.520 1.850 ;
        RECT  8.495 1.590 8.920 1.750 ;
        RECT  8.515 2.165 8.775 2.425 ;
        RECT  8.405 2.615 8.565 3.105 ;
        RECT  7.445 2.265 8.515 2.425 ;
        RECT  8.335 1.145 8.495 1.750 ;
        RECT  7.135 2.945 8.405 3.105 ;
        RECT  6.995 1.145 8.335 1.305 ;
        RECT  6.995 2.605 8.225 2.765 ;
        RECT  7.735 0.595 7.785 0.915 ;
        RECT  7.525 0.595 7.735 0.965 ;
        RECT  5.480 0.805 7.525 0.965 ;
        RECT  7.285 1.680 7.445 2.425 ;
        RECT  7.185 1.680 7.285 1.940 ;
        RECT  6.875 2.945 7.135 3.205 ;
        RECT  6.835 1.145 6.995 2.765 ;
        RECT  6.165 2.945 6.875 3.105 ;
        RECT  6.045 1.195 6.835 1.355 ;
        RECT  6.705 2.505 6.835 2.765 ;
        RECT  5.625 2.605 6.705 2.765 ;
        RECT  6.495 1.740 6.655 2.250 ;
        RECT  5.295 1.740 6.495 1.900 ;
        RECT  6.005 2.945 6.165 3.220 ;
        RECT  5.785 1.145 6.045 1.405 ;
        RECT  4.960 3.060 6.005 3.220 ;
        RECT  5.365 2.275 5.625 2.875 ;
        RECT  5.320 0.805 5.480 1.240 ;
        RECT  4.425 1.080 5.320 1.240 ;
        RECT  5.140 1.525 5.295 1.900 ;
        RECT  4.880 0.535 5.140 0.795 ;
        RECT  5.135 1.425 5.140 1.900 ;
        RECT  4.880 1.425 5.135 1.685 ;
        RECT  4.800 2.945 4.960 3.220 ;
        RECT  3.090 0.585 4.880 0.745 ;
        RECT  4.425 1.985 4.855 2.245 ;
        RECT  0.810 2.945 4.800 3.105 ;
        RECT  4.265 1.080 4.425 2.665 ;
        RECT  3.475 1.080 4.265 1.240 ;
        RECT  4.080 2.505 4.265 2.665 ;
        RECT  3.820 2.505 4.080 2.765 ;
        RECT  2.690 2.605 3.820 2.765 ;
        RECT  3.215 1.030 3.475 1.290 ;
        RECT  3.030 2.265 3.130 2.425 ;
        RECT  3.030 0.520 3.090 0.780 ;
        RECT  2.870 0.520 3.030 2.425 ;
        RECT  2.830 0.520 2.870 0.780 ;
        RECT  2.530 1.685 2.690 2.765 ;
        RECT  2.410 1.685 2.530 1.845 ;
        RECT  2.150 1.585 2.410 1.845 ;
        RECT  1.960 2.165 2.220 2.765 ;
        RECT  1.935 0.430 2.095 0.745 ;
        RECT  1.270 2.170 1.960 2.330 ;
        RECT  0.470 0.585 1.935 0.745 ;
        RECT  1.300 0.930 1.560 1.190 ;
        RECT  0.810 1.030 1.300 1.190 ;
        RECT  1.010 1.955 1.270 2.330 ;
        RECT  0.650 1.030 0.810 3.105 ;
        RECT  0.310 0.585 0.470 2.855 ;
        RECT  0.210 0.900 0.310 1.160 ;
        RECT  0.210 2.595 0.310 2.855 ;
    END
END DFFSHQX8

MACRO DFFSHQX4
    CLASS CORE ;
    FOREIGN DFFSHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.640 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.660 1.700 8.155 2.085 ;
        END
        ANTENNAGATEAREA     0.3510 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.795 0.600 15.055 3.060 ;
        END
        ANTENNADIFFAREA     0.8132 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.620 3.715 1.990 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.495 1.715 1.990 ;
        RECT  1.350 1.495 1.505 1.755 ;
        END
        ANTENNAGATEAREA     0.4563 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.515 -0.250 15.640 0.250 ;
        RECT  15.255 -0.250 15.515 1.095 ;
        RECT  14.440 -0.250 15.255 0.250 ;
        RECT  14.180 -0.250 14.440 0.405 ;
        RECT  12.300 -0.250 14.180 0.250 ;
        RECT  12.660 1.000 12.920 1.260 ;
        RECT  12.300 1.000 12.660 1.160 ;
        RECT  12.140 -0.250 12.300 1.160 ;
        RECT  9.980 -0.250 12.140 0.250 ;
        RECT  9.720 -0.250 9.980 0.575 ;
        RECT  8.895 -0.250 9.720 0.250 ;
        RECT  8.635 -0.250 8.895 0.575 ;
        RECT  8.325 -0.250 8.635 0.250 ;
        RECT  8.065 -0.250 8.325 0.575 ;
        RECT  7.225 -0.250 8.065 0.250 ;
        RECT  6.965 -0.250 7.225 0.625 ;
        RECT  4.030 -0.250 6.965 0.250 ;
        RECT  3.770 -0.250 4.030 0.405 ;
        RECT  2.535 -0.250 3.770 0.250 ;
        RECT  2.275 -0.250 2.535 1.065 ;
        RECT  1.020 -0.250 2.275 0.250 ;
        RECT  0.760 -0.250 1.020 0.405 ;
        RECT  0.000 -0.250 0.760 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.515 3.440 15.640 3.940 ;
        RECT  15.255 2.275 15.515 3.940 ;
        RECT  14.340 3.440 15.255 3.940 ;
        RECT  14.080 3.285 14.340 3.940 ;
        RECT  11.890 3.440 14.080 3.940 ;
        RECT  11.630 3.285 11.890 3.940 ;
        RECT  9.285 3.440 11.630 3.940 ;
        RECT  9.025 2.955 9.285 3.940 ;
        RECT  7.675 3.440 9.025 3.940 ;
        RECT  7.415 3.285 7.675 3.940 ;
        RECT  6.605 3.440 7.415 3.940 ;
        RECT  6.345 3.285 6.605 3.940 ;
        RECT  4.620 3.440 6.345 3.940 ;
        RECT  4.360 3.285 4.620 3.940 ;
        RECT  3.530 3.440 4.360 3.940 ;
        RECT  3.270 3.285 3.530 3.940 ;
        RECT  1.670 3.440 3.270 3.940 ;
        RECT  1.410 3.285 1.670 3.940 ;
        RECT  0.000 3.440 1.410 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.400 0.590 14.560 3.105 ;
        RECT  14.000 0.590 14.400 0.750 ;
        RECT  13.520 2.945 14.400 3.105 ;
        RECT  14.060 1.640 14.220 2.750 ;
        RECT  13.780 1.640 14.060 1.900 ;
        RECT  13.080 2.590 14.060 2.750 ;
        RECT  13.840 0.470 14.000 0.750 ;
        RECT  13.440 2.245 13.880 2.405 ;
        RECT  12.660 0.470 13.840 0.630 ;
        RECT  13.660 0.930 13.780 1.900 ;
        RECT  13.620 0.810 13.660 1.900 ;
        RECT  13.400 0.810 13.620 1.090 ;
        RECT  13.360 2.945 13.520 3.260 ;
        RECT  13.280 1.270 13.440 2.405 ;
        RECT  12.790 3.100 13.360 3.260 ;
        RECT  12.305 1.765 13.280 1.925 ;
        RECT  12.920 2.590 13.080 2.865 ;
        RECT  11.625 2.705 12.920 2.865 ;
        RECT  12.480 2.265 12.740 2.525 ;
        RECT  11.965 2.265 12.480 2.425 ;
        RECT  12.145 1.765 12.305 2.045 ;
        RECT  11.900 1.555 11.965 2.425 ;
        RECT  11.805 0.470 11.900 2.425 ;
        RECT  11.740 0.470 11.805 1.715 ;
        RECT  10.320 0.470 11.740 0.630 ;
        RECT  11.560 1.905 11.625 2.865 ;
        RECT  11.465 0.810 11.560 2.865 ;
        RECT  11.400 0.810 11.465 2.065 ;
        RECT  10.660 0.810 11.400 0.970 ;
        RECT  10.825 1.905 11.400 2.065 ;
        RECT  11.125 2.255 11.285 3.220 ;
        RECT  10.385 3.060 11.125 3.220 ;
        RECT  11.000 1.155 11.100 1.315 ;
        RECT  10.840 1.155 11.000 1.725 ;
        RECT  10.385 1.565 10.840 1.725 ;
        RECT  10.615 1.905 10.825 2.875 ;
        RECT  10.500 0.810 10.660 1.315 ;
        RECT  10.565 2.275 10.615 2.875 ;
        RECT  10.205 1.155 10.500 1.315 ;
        RECT  10.225 1.565 10.385 3.220 ;
        RECT  10.205 0.470 10.320 0.915 ;
        RECT  9.870 2.165 10.225 2.425 ;
        RECT  10.160 0.470 10.205 0.945 ;
        RECT  9.945 0.755 10.160 0.945 ;
        RECT  9.845 2.615 10.005 3.215 ;
        RECT  7.785 0.755 9.945 0.915 ;
        RECT  9.710 1.115 9.870 2.425 ;
        RECT  8.565 2.615 9.845 2.775 ;
        RECT  9.175 1.115 9.710 1.275 ;
        RECT  9.535 2.165 9.710 2.425 ;
        RECT  8.775 2.265 9.535 2.425 ;
        RECT  8.895 1.590 9.495 1.850 ;
        RECT  8.495 1.590 8.895 1.750 ;
        RECT  8.515 2.165 8.775 2.425 ;
        RECT  8.405 2.615 8.565 3.105 ;
        RECT  7.445 2.265 8.515 2.425 ;
        RECT  8.335 1.145 8.495 1.750 ;
        RECT  7.135 2.945 8.405 3.105 ;
        RECT  6.995 1.145 8.335 1.305 ;
        RECT  6.995 2.605 8.225 2.765 ;
        RECT  7.735 0.475 7.785 0.915 ;
        RECT  7.525 0.475 7.735 0.965 ;
        RECT  5.480 0.805 7.525 0.965 ;
        RECT  7.285 1.680 7.445 2.425 ;
        RECT  7.185 1.680 7.285 1.940 ;
        RECT  6.875 2.945 7.135 3.205 ;
        RECT  6.835 1.145 6.995 2.765 ;
        RECT  6.165 2.945 6.875 3.105 ;
        RECT  6.045 1.195 6.835 1.355 ;
        RECT  6.705 2.505 6.835 2.765 ;
        RECT  5.625 2.605 6.705 2.765 ;
        RECT  6.495 1.740 6.655 2.250 ;
        RECT  5.295 1.740 6.495 1.900 ;
        RECT  6.005 2.945 6.165 3.220 ;
        RECT  5.785 1.145 6.045 1.405 ;
        RECT  4.960 3.060 6.005 3.220 ;
        RECT  5.365 2.275 5.625 2.875 ;
        RECT  5.320 0.805 5.480 1.240 ;
        RECT  4.425 1.080 5.320 1.240 ;
        RECT  5.140 1.525 5.295 1.900 ;
        RECT  4.880 0.535 5.140 0.795 ;
        RECT  5.135 1.425 5.140 1.900 ;
        RECT  4.880 1.425 5.135 1.685 ;
        RECT  4.800 2.945 4.960 3.220 ;
        RECT  3.090 0.585 4.880 0.745 ;
        RECT  4.425 1.985 4.855 2.245 ;
        RECT  0.830 2.945 4.800 3.105 ;
        RECT  4.265 1.080 4.425 2.665 ;
        RECT  3.475 1.080 4.265 1.240 ;
        RECT  4.080 2.505 4.265 2.665 ;
        RECT  3.820 2.505 4.080 2.765 ;
        RECT  2.690 2.605 3.820 2.765 ;
        RECT  3.215 1.030 3.475 1.290 ;
        RECT  3.030 2.265 3.130 2.425 ;
        RECT  3.030 0.520 3.090 0.780 ;
        RECT  2.870 0.520 3.030 2.425 ;
        RECT  2.830 0.520 2.870 0.780 ;
        RECT  2.530 1.685 2.690 2.765 ;
        RECT  2.390 1.685 2.530 1.845 ;
        RECT  2.130 1.585 2.390 1.845 ;
        RECT  1.960 2.165 2.220 2.765 ;
        RECT  1.835 0.535 2.095 0.795 ;
        RECT  1.270 2.170 1.960 2.330 ;
        RECT  0.470 0.585 1.835 0.745 ;
        RECT  1.300 0.935 1.560 1.195 ;
        RECT  0.830 1.035 1.300 1.195 ;
        RECT  1.010 1.955 1.270 2.330 ;
        RECT  0.670 1.035 0.830 3.105 ;
        RECT  0.310 0.585 0.470 2.865 ;
        RECT  0.210 0.900 0.310 1.160 ;
        RECT  0.210 2.605 0.310 2.865 ;
    END
END DFFSHQX4

MACRO DFFSHQX2
    CLASS CORE ;
    FOREIGN DFFSHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.240 1.575 6.500 2.075 ;
        RECT  6.065 1.630 6.240 2.075 ;
        END
        ANTENNAGATEAREA     0.2054 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.395 0.600 11.550 1.355 ;
        RECT  11.290 0.600 11.395 2.600 ;
        RECT  11.235 0.695 11.290 2.600 ;
        RECT  11.165 1.515 11.235 2.600 ;
        RECT  11.135 2.000 11.165 2.600 ;
        END
        ANTENNADIFFAREA     0.5668 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 1.700 3.095 2.005 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.470 0.950 1.990 ;
        END
        ANTENNAGATEAREA     0.2626 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.010 -0.250 11.960 0.250 ;
        RECT  10.750 -0.250 11.010 1.050 ;
        RECT  8.535 -0.250 10.750 0.250 ;
        RECT  8.275 -0.250 8.535 0.405 ;
        RECT  6.745 -0.250 8.275 0.250 ;
        RECT  6.485 -0.250 6.745 0.405 ;
        RECT  6.120 -0.250 6.485 0.250 ;
        RECT  5.960 -0.250 6.120 0.655 ;
        RECT  3.650 -0.250 5.960 0.250 ;
        RECT  3.390 -0.250 3.650 0.405 ;
        RECT  2.675 -0.250 3.390 0.250 ;
        RECT  2.415 -0.250 2.675 0.405 ;
        RECT  0.930 -0.250 2.415 0.250 ;
        RECT  0.670 -0.250 0.930 0.405 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.795 3.440 11.960 3.940 ;
        RECT  11.195 3.060 11.795 3.940 ;
        RECT  8.555 3.440 11.195 3.940 ;
        RECT  8.295 2.965 8.555 3.940 ;
        RECT  7.005 3.440 8.295 3.940 ;
        RECT  6.745 3.115 7.005 3.940 ;
        RECT  5.405 3.440 6.745 3.940 ;
        RECT  5.145 3.285 5.405 3.940 ;
        RECT  3.755 3.440 5.145 3.940 ;
        RECT  3.495 3.285 3.755 3.940 ;
        RECT  2.705 3.440 3.495 3.940 ;
        RECT  2.445 3.285 2.705 3.940 ;
        RECT  0.920 3.440 2.445 3.940 ;
        RECT  0.660 2.890 0.920 3.940 ;
        RECT  0.000 3.440 0.660 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.745 1.230 10.905 3.165 ;
        RECT  10.510 1.230 10.745 1.390 ;
        RECT  10.395 3.005 10.745 3.165 ;
        RECT  10.355 1.570 10.515 2.790 ;
        RECT  10.350 0.430 10.510 1.390 ;
        RECT  9.720 3.005 10.395 3.235 ;
        RECT  10.255 1.570 10.355 1.830 ;
        RECT  9.120 2.630 10.355 2.790 ;
        RECT  9.730 0.430 10.350 0.590 ;
        RECT  10.170 1.570 10.255 1.730 ;
        RECT  10.010 0.770 10.170 1.730 ;
        RECT  10.010 2.010 10.170 2.270 ;
        RECT  9.910 0.770 10.010 0.930 ;
        RECT  9.830 2.010 10.010 2.170 ;
        RECT  9.670 1.325 9.830 2.170 ;
        RECT  9.570 0.430 9.730 0.645 ;
        RECT  9.590 1.325 9.670 1.485 ;
        RECT  9.330 1.035 9.590 1.485 ;
        RECT  9.115 0.485 9.570 0.645 ;
        RECT  9.305 1.665 9.465 2.450 ;
        RECT  8.905 1.325 9.330 1.485 ;
        RECT  8.395 1.665 9.305 1.825 ;
        RECT  8.960 2.045 9.120 2.790 ;
        RECT  8.855 0.485 9.115 0.785 ;
        RECT  8.055 2.045 8.960 2.205 ;
        RECT  8.645 1.225 8.905 1.485 ;
        RECT  8.305 2.385 8.565 2.645 ;
        RECT  8.235 0.585 8.395 1.825 ;
        RECT  7.545 2.435 8.305 2.595 ;
        RECT  8.055 0.585 8.235 0.745 ;
        RECT  7.795 0.430 8.055 0.745 ;
        RECT  7.955 1.995 8.055 2.255 ;
        RECT  7.795 0.925 7.955 2.255 ;
        RECT  7.545 2.775 7.805 3.215 ;
        RECT  6.775 0.585 7.795 0.745 ;
        RECT  7.535 0.925 7.795 1.185 ;
        RECT  7.355 2.310 7.545 2.595 ;
        RECT  6.295 2.775 7.545 2.935 ;
        RECT  7.195 0.925 7.355 2.595 ;
        RECT  7.025 0.925 7.195 1.185 ;
        RECT  6.465 2.435 7.195 2.595 ;
        RECT  6.840 1.400 7.015 2.000 ;
        RECT  6.755 1.175 6.840 2.000 ;
        RECT  6.615 0.585 6.775 0.995 ;
        RECT  6.680 1.175 6.755 1.560 ;
        RECT  6.005 1.175 6.680 1.335 ;
        RECT  5.750 0.835 6.615 0.995 ;
        RECT  6.205 2.265 6.465 2.595 ;
        RECT  6.135 2.775 6.295 3.105 ;
        RECT  5.255 2.265 6.205 2.425 ;
        RECT  4.865 2.945 6.135 3.105 ;
        RECT  5.845 1.175 6.005 1.415 ;
        RECT  4.850 2.605 5.955 2.765 ;
        RECT  4.850 1.255 5.845 1.415 ;
        RECT  5.665 0.475 5.750 0.995 ;
        RECT  5.500 0.475 5.665 1.075 ;
        RECT  4.510 0.915 5.500 1.075 ;
        RECT  5.060 0.475 5.320 0.735 ;
        RECT  5.095 1.710 5.255 2.425 ;
        RECT  4.165 0.475 5.060 0.635 ;
        RECT  4.605 2.945 4.865 3.205 ;
        RECT  4.690 1.255 4.850 2.765 ;
        RECT  4.395 2.325 4.690 2.765 ;
        RECT  4.215 2.945 4.605 3.105 ;
        RECT  4.350 0.915 4.510 1.425 ;
        RECT  4.215 1.605 4.410 1.865 ;
        RECT  3.875 1.265 4.350 1.425 ;
        RECT  4.055 1.605 4.215 3.105 ;
        RECT  4.005 0.475 4.165 1.085 ;
        RECT  1.290 2.945 4.055 3.105 ;
        RECT  2.205 0.925 4.005 1.085 ;
        RECT  3.715 1.265 3.875 2.765 ;
        RECT  2.925 1.265 3.715 1.425 ;
        RECT  3.215 2.605 3.715 2.765 ;
        RECT  2.955 2.335 3.215 2.765 ;
        RECT  3.000 0.435 3.160 0.745 ;
        RECT  0.405 0.585 3.000 0.745 ;
        RECT  1.730 2.605 2.955 2.765 ;
        RECT  2.205 2.165 2.305 2.425 ;
        RECT  2.045 0.925 2.205 2.425 ;
        RECT  1.845 0.925 2.045 1.185 ;
        RECT  1.570 1.655 1.730 2.765 ;
        RECT  1.470 1.655 1.570 1.915 ;
        RECT  1.290 1.035 1.500 1.295 ;
        RECT  1.130 1.035 1.290 3.105 ;
        RECT  0.405 2.185 0.520 2.445 ;
        RECT  0.245 0.585 0.405 2.445 ;
        RECT  0.125 1.035 0.245 1.295 ;
    END
END DFFSHQX2

MACRO DFFSHQX1
    CLASS CORE ;
    FOREIGN DFFSHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 1.700 6.775 1.990 ;
        RECT  5.945 1.700 6.565 1.865 ;
        RECT  5.785 1.555 5.945 1.865 ;
        END
        ANTENNAGATEAREA     0.1352 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.535 1.990 9.670 2.250 ;
        RECT  9.510 1.515 9.535 2.250 ;
        RECT  9.485 1.515 9.510 2.150 ;
        RECT  9.325 0.930 9.485 2.150 ;
        RECT  9.185 0.930 9.325 1.190 ;
        END
        ANTENNADIFFAREA     0.3861 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 1.700 2.185 2.240 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.540 0.840 1.990 ;
        RECT  0.495 1.545 0.585 1.805 ;
        END
        ANTENNAGATEAREA     0.1560 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.215 -0.250 10.580 0.250 ;
        RECT  9.955 -0.250 10.215 0.405 ;
        RECT  8.095 -0.250 9.955 0.250 ;
        RECT  7.835 -0.250 8.095 0.405 ;
        RECT  6.325 -0.250 7.835 0.250 ;
        RECT  6.065 -0.250 6.325 0.405 ;
        RECT  5.750 -0.250 6.065 0.250 ;
        RECT  5.490 -0.250 5.750 0.655 ;
        RECT  3.285 -0.250 5.490 0.250 ;
        RECT  3.025 -0.250 3.285 0.405 ;
        RECT  1.305 -0.250 3.025 0.250 ;
        RECT  0.705 -0.250 1.305 0.405 ;
        RECT  0.000 -0.250 0.705 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.980 3.440 10.580 3.940 ;
        RECT  9.040 3.115 9.980 3.940 ;
        RECT  6.060 3.440 9.040 3.940 ;
        RECT  5.800 3.115 6.060 3.940 ;
        RECT  5.100 3.440 5.800 3.940 ;
        RECT  4.840 3.285 5.100 3.940 ;
        RECT  3.295 3.440 4.840 3.940 ;
        RECT  3.035 3.285 3.295 3.940 ;
        RECT  2.195 3.440 3.035 3.940 ;
        RECT  1.935 3.285 2.195 3.940 ;
        RECT  0.810 3.440 1.935 3.940 ;
        RECT  0.550 2.890 0.810 3.940 ;
        RECT  0.000 3.440 0.550 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.375 0.585 10.485 1.500 ;
        RECT  10.350 0.585 10.375 1.600 ;
        RECT  10.325 0.585 10.350 2.935 ;
        RECT  9.475 0.585 10.325 0.745 ;
        RECT  10.190 1.340 10.325 2.935 ;
        RECT  8.625 2.775 10.190 2.935 ;
        RECT  10.010 1.000 10.145 1.160 ;
        RECT  9.850 1.000 10.010 2.590 ;
        RECT  9.060 2.430 9.850 2.590 ;
        RECT  9.310 0.430 9.475 0.745 ;
        RECT  9.215 0.430 9.310 0.590 ;
        RECT  9.060 1.460 9.105 1.720 ;
        RECT  9.005 1.460 9.060 2.590 ;
        RECT  8.900 0.640 9.005 2.590 ;
        RECT  8.845 0.640 8.900 1.720 ;
        RECT  8.270 2.345 8.900 2.505 ;
        RECT  7.505 0.640 8.845 0.800 ;
        RECT  8.530 1.905 8.720 2.165 ;
        RECT  8.465 2.775 8.625 3.165 ;
        RECT  8.370 0.980 8.530 2.165 ;
        RECT  7.600 3.005 8.465 3.165 ;
        RECT  8.270 0.980 8.370 1.240 ;
        RECT  7.870 1.725 8.370 1.985 ;
        RECT  8.110 2.345 8.270 2.710 ;
        RECT  7.115 2.550 8.110 2.710 ;
        RECT  7.345 0.465 7.505 0.800 ;
        RECT  7.455 1.570 7.460 2.295 ;
        RECT  7.300 1.005 7.455 2.295 ;
        RECT  6.605 3.005 7.375 3.165 ;
        RECT  7.295 1.005 7.300 1.730 ;
        RECT  7.165 1.005 7.295 1.165 ;
        RECT  7.005 0.585 7.165 1.165 ;
        RECT  6.955 1.360 7.115 2.330 ;
        RECT  6.855 2.550 7.115 2.810 ;
        RECT  6.900 0.585 7.005 0.745 ;
        RECT  6.825 1.360 6.955 1.520 ;
        RECT  6.600 2.170 6.955 2.330 ;
        RECT  6.640 0.450 6.900 0.745 ;
        RECT  6.665 0.925 6.825 1.520 ;
        RECT  6.470 0.925 6.665 1.085 ;
        RECT  6.270 0.585 6.640 0.745 ;
        RECT  6.445 2.770 6.605 3.165 ;
        RECT  6.340 2.170 6.600 2.590 ;
        RECT  6.285 1.360 6.475 1.520 ;
        RECT  5.285 2.770 6.445 2.935 ;
        RECT  6.030 2.170 6.340 2.330 ;
        RECT  6.125 1.215 6.285 1.520 ;
        RECT  6.110 0.585 6.270 0.995 ;
        RECT  5.550 1.215 6.125 1.375 ;
        RECT  5.205 0.835 6.110 0.995 ;
        RECT  5.870 2.045 6.030 2.330 ;
        RECT  5.515 2.045 5.870 2.205 ;
        RECT  4.705 2.385 5.690 2.545 ;
        RECT  5.390 1.215 5.550 1.445 ;
        RECT  5.355 1.625 5.515 2.205 ;
        RECT  4.705 1.285 5.390 1.445 ;
        RECT  5.255 1.625 5.355 1.785 ;
        RECT  5.120 2.770 5.285 3.105 ;
        RECT  5.105 0.475 5.205 0.995 ;
        RECT  4.595 2.945 5.120 3.105 ;
        RECT  4.945 0.475 5.105 1.105 ;
        RECT  2.980 0.930 4.945 1.105 ;
        RECT  4.460 0.475 4.720 0.745 ;
        RECT  4.545 1.285 4.705 2.545 ;
        RECT  4.335 2.895 4.595 3.155 ;
        RECT  4.315 1.285 4.545 1.445 ;
        RECT  4.145 2.275 4.545 2.545 ;
        RECT  2.415 0.585 4.460 0.745 ;
        RECT  3.965 2.945 4.335 3.105 ;
        RECT  3.805 1.585 3.965 3.105 ;
        RECT  3.545 1.585 3.805 1.745 ;
        RECT  1.685 2.945 3.805 3.105 ;
        RECT  2.980 2.015 3.615 2.275 ;
        RECT  2.820 0.930 2.980 2.765 ;
        RECT  2.595 0.930 2.820 1.090 ;
        RECT  1.625 2.605 2.820 2.765 ;
        RECT  2.535 1.805 2.635 2.065 ;
        RECT  2.415 1.345 2.535 2.065 ;
        RECT  2.375 0.585 2.415 2.065 ;
        RECT  2.255 0.585 2.375 1.505 ;
        RECT  1.865 0.585 2.255 0.845 ;
        RECT  1.915 1.025 2.075 1.285 ;
        RECT  1.685 1.025 1.915 1.185 ;
        RECT  1.525 0.690 1.685 1.185 ;
        RECT  1.425 2.945 1.685 3.215 ;
        RECT  1.465 1.815 1.625 2.765 ;
        RECT  0.385 0.690 1.525 0.850 ;
        RECT  1.365 1.815 1.465 2.075 ;
        RECT  1.185 2.945 1.425 3.105 ;
        RECT  1.185 1.035 1.345 1.295 ;
        RECT  1.025 1.135 1.185 3.105 ;
        RECT  0.285 0.690 0.385 1.295 ;
        RECT  0.285 2.185 0.385 2.445 ;
        RECT  0.225 0.690 0.285 2.445 ;
        RECT  0.125 1.035 0.225 2.445 ;
    END
END DFFSHQX1

MACRO DFFRHQX8
    CLASS CORE ;
    FOREIGN DFFRHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.280 1.885 10.440 2.145 ;
        RECT  8.130 1.985 10.280 2.145 ;
        RECT  8.155 1.275 8.190 1.535 ;
        RECT  8.130 1.275 8.155 1.700 ;
        RECT  8.105 1.275 8.130 2.145 ;
        RECT  8.030 1.275 8.105 2.170 ;
        RECT  7.945 1.290 8.030 2.170 ;
        RECT  6.940 1.295 7.945 1.455 ;
        RECT  7.665 2.010 7.945 2.170 ;
        RECT  6.680 1.295 6.940 1.485 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.000 1.515 14.135 1.765 ;
        RECT  13.740 0.695 14.000 3.055 ;
        RECT  13.215 1.300 13.740 1.705 ;
        RECT  12.980 1.300 13.215 2.400 ;
        RECT  12.720 0.695 12.980 3.055 ;
        RECT  12.545 1.515 12.720 2.585 ;
        END
        ANTENNADIFFAREA     1.6264 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.490 2.360 1.990 ;
        END
        ANTENNAGATEAREA     0.1534 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.445 0.425 1.990 ;
        END
        ANTENNAGATEAREA     0.3744 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.510 -0.250 14.720 0.250 ;
        RECT  14.250 -0.250 14.510 1.095 ;
        RECT  13.490 -0.250 14.250 0.250 ;
        RECT  13.230 -0.250 13.490 1.120 ;
        RECT  12.440 -0.250 13.230 0.250 ;
        RECT  12.180 -0.250 12.440 0.840 ;
        RECT  11.230 -0.250 12.180 0.250 ;
        RECT  10.970 -0.250 11.230 0.405 ;
        RECT  8.560 -0.250 10.970 0.250 ;
        RECT  8.300 -0.250 8.560 0.405 ;
        RECT  6.695 -0.250 8.300 0.250 ;
        RECT  6.435 -0.250 6.695 0.405 ;
        RECT  5.590 -0.250 6.435 0.250 ;
        RECT  5.330 -0.250 5.590 0.405 ;
        RECT  3.830 -0.250 5.330 0.250 ;
        RECT  3.670 -0.250 3.830 0.935 ;
        RECT  2.470 -0.250 3.670 0.250 ;
        RECT  2.210 -0.250 2.470 0.870 ;
        RECT  0.945 -0.250 2.210 0.250 ;
        RECT  0.685 -0.250 0.945 0.405 ;
        RECT  0.000 -0.250 0.685 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.510 3.440 14.720 3.940 ;
        RECT  14.250 2.275 14.510 3.940 ;
        RECT  13.490 3.440 14.250 3.940 ;
        RECT  13.230 2.615 13.490 3.940 ;
        RECT  12.280 3.440 13.230 3.940 ;
        RECT  12.020 2.955 12.280 3.940 ;
        RECT  10.870 3.440 12.020 3.940 ;
        RECT  10.610 3.065 10.870 3.940 ;
        RECT  7.500 3.440 10.610 3.940 ;
        RECT  7.240 3.285 7.500 3.940 ;
        RECT  6.400 3.440 7.240 3.940 ;
        RECT  6.140 3.285 6.400 3.940 ;
        RECT  5.145 3.440 6.140 3.940 ;
        RECT  4.885 3.285 5.145 3.940 ;
        RECT  3.410 3.440 4.885 3.940 ;
        RECT  3.150 3.285 3.410 3.940 ;
        RECT  2.460 3.440 3.150 3.940 ;
        RECT  2.200 3.285 2.460 3.940 ;
        RECT  0.765 3.440 2.200 3.940 ;
        RECT  0.505 2.955 0.765 3.940 ;
        RECT  0.000 3.440 0.505 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.350 1.545 12.355 1.805 ;
        RECT  12.190 1.545 12.350 2.505 ;
        RECT  12.095 1.545 12.190 1.805 ;
        RECT  12.170 2.345 12.190 2.505 ;
        RECT  12.010 2.345 12.170 2.775 ;
        RECT  11.800 2.005 12.010 2.165 ;
        RECT  11.675 2.615 12.010 2.775 ;
        RECT  11.640 1.035 11.800 2.165 ;
        RECT  11.415 2.615 11.675 2.880 ;
        RECT  11.300 0.585 11.460 2.435 ;
        RECT  11.120 2.665 11.415 2.825 ;
        RECT  9.640 0.585 11.300 0.745 ;
        RECT  10.960 0.925 11.120 2.825 ;
        RECT  8.870 0.925 10.960 1.085 ;
        RECT  9.655 2.665 10.960 2.825 ;
        RECT  10.620 1.365 10.780 2.485 ;
        RECT  9.500 1.365 10.620 1.525 ;
        RECT  9.145 2.325 10.620 2.485 ;
        RECT  10.165 3.005 10.425 3.220 ;
        RECT  7.870 3.060 10.165 3.220 ;
        RECT  9.425 2.665 9.655 2.880 ;
        RECT  9.040 0.440 9.640 0.745 ;
        RECT  9.240 1.265 9.500 1.525 ;
        RECT  8.375 2.720 9.425 2.880 ;
        RECT  8.530 1.365 9.240 1.525 ;
        RECT  8.980 2.325 9.145 2.540 ;
        RECT  6.150 0.585 9.040 0.745 ;
        RECT  8.125 2.380 8.980 2.540 ;
        RECT  8.710 0.925 8.870 1.185 ;
        RECT  8.370 0.925 8.530 1.525 ;
        RECT  7.330 0.925 8.370 1.085 ;
        RECT  7.865 2.380 8.125 2.715 ;
        RECT  7.710 2.945 7.870 3.220 ;
        RECT  6.950 2.380 7.865 2.540 ;
        RECT  5.705 2.945 7.710 3.105 ;
        RECT  7.185 1.635 7.445 1.825 ;
        RECT  6.470 1.665 7.185 1.825 ;
        RECT  6.690 2.165 6.950 2.765 ;
        RECT  6.130 2.165 6.690 2.325 ;
        RECT  6.310 1.085 6.470 1.825 ;
        RECT  5.720 1.085 6.310 1.245 ;
        RECT  5.890 0.510 6.150 0.905 ;
        RECT  5.970 1.430 6.130 2.325 ;
        RECT  4.180 0.745 5.890 0.905 ;
        RECT  5.560 1.085 5.720 2.275 ;
        RECT  5.545 2.560 5.705 3.105 ;
        RECT  4.470 1.085 5.560 1.245 ;
        RECT  5.505 2.115 5.560 2.275 ;
        RECT  5.445 2.560 5.545 3.055 ;
        RECT  5.245 2.115 5.505 2.380 ;
        RECT  5.440 2.610 5.445 3.055 ;
        RECT  3.835 2.895 5.440 3.055 ;
        RECT  5.280 1.460 5.380 1.620 ;
        RECT  5.120 1.460 5.280 1.870 ;
        RECT  4.275 2.115 5.245 2.275 ;
        RECT  4.080 1.710 5.120 1.870 ;
        RECT  4.015 2.115 4.275 2.715 ;
        RECT  4.020 0.745 4.180 1.275 ;
        RECT  3.835 1.455 4.080 1.870 ;
        RECT  3.440 1.115 4.020 1.275 ;
        RECT  3.820 1.455 3.835 3.055 ;
        RECT  3.675 1.710 3.820 3.055 ;
        RECT  1.105 2.895 3.675 3.055 ;
        RECT  3.300 0.455 3.460 0.715 ;
        RECT  3.280 1.115 3.440 2.255 ;
        RECT  2.810 0.555 3.300 0.715 ;
        RECT  3.250 1.115 3.280 1.275 ;
        RECT  3.010 2.095 3.280 2.255 ;
        RECT  3.040 0.895 3.250 1.275 ;
        RECT  2.990 0.895 3.040 1.155 ;
        RECT  2.750 2.095 3.010 2.715 ;
        RECT  2.650 0.555 2.810 1.295 ;
        RECT  1.445 2.555 2.750 2.715 ;
        RECT  1.930 1.135 2.650 1.295 ;
        RECT  1.785 2.215 2.060 2.375 ;
        RECT  1.785 0.950 1.930 1.295 ;
        RECT  1.740 0.480 1.790 0.740 ;
        RECT  1.670 0.950 1.785 2.375 ;
        RECT  1.530 0.480 1.740 0.745 ;
        RECT  1.625 1.135 1.670 2.375 ;
        RECT  0.765 0.585 1.530 0.745 ;
        RECT  1.285 1.580 1.445 2.715 ;
        RECT  1.105 1.035 1.345 1.295 ;
        RECT  0.945 1.035 1.105 3.055 ;
        RECT  0.605 0.585 0.765 2.345 ;
        RECT  0.135 0.905 0.605 1.165 ;
        RECT  0.395 2.185 0.605 2.345 ;
        RECT  0.135 2.185 0.395 2.445 ;
    END
END DFFRHQX8

MACRO DFFRHQX4
    CLASS CORE ;
    FOREIGN DFFRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.340 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.905 1.705 10.065 2.045 ;
        RECT  8.055 1.705 9.905 1.865 ;
        RECT  7.895 1.280 8.055 1.865 ;
        RECT  6.775 1.280 7.895 1.440 ;
        RECT  6.565 1.280 6.775 1.580 ;
        END
        ANTENNAGATEAREA     0.3874 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.425 0.590 12.685 1.190 ;
        RECT  12.295 2.140 12.430 3.080 ;
        RECT  12.295 0.880 12.425 1.190 ;
        RECT  12.270 0.880 12.295 3.080 ;
        RECT  12.170 0.990 12.270 3.080 ;
        RECT  12.095 0.990 12.170 2.585 ;
        RECT  12.085 1.170 12.095 2.585 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.700 2.635 1.990 ;
        RECT  2.165 1.700 2.425 1.860 ;
        RECT  2.005 1.585 2.165 1.860 ;
        END
        ANTENNAGATEAREA     0.1534 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.420 0.795 1.990 ;
        RECT  0.470 1.420 0.585 1.905 ;
        END
        ANTENNAGATEAREA     0.3744 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.195 -0.250 13.340 0.250 ;
        RECT  12.935 -0.250 13.195 1.165 ;
        RECT  12.135 -0.250 12.935 0.250 ;
        RECT  11.875 -0.250 12.135 0.405 ;
        RECT  10.915 -0.250 11.875 0.250 ;
        RECT  10.655 -0.250 10.915 0.405 ;
        RECT  8.315 -0.250 10.655 0.250 ;
        RECT  8.055 -0.250 8.315 0.405 ;
        RECT  6.555 -0.250 8.055 0.250 ;
        RECT  6.295 -0.250 6.555 0.565 ;
        RECT  5.455 -0.250 6.295 0.250 ;
        RECT  5.195 -0.250 5.455 0.405 ;
        RECT  3.445 -0.250 5.195 0.250 ;
        RECT  3.185 -0.250 3.445 0.405 ;
        RECT  2.335 -0.250 3.185 0.250 ;
        RECT  2.175 -0.250 2.335 0.955 ;
        RECT  0.785 -0.250 2.175 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.940 3.440 13.340 3.940 ;
        RECT  12.680 2.230 12.940 3.940 ;
        RECT  11.685 3.440 12.680 3.940 ;
        RECT  11.425 2.935 11.685 3.940 ;
        RECT  10.225 3.440 11.425 3.940 ;
        RECT  9.965 3.065 10.225 3.940 ;
        RECT  7.530 3.440 9.965 3.940 ;
        RECT  7.270 3.285 7.530 3.940 ;
        RECT  6.310 3.440 7.270 3.940 ;
        RECT  6.050 3.285 6.310 3.940 ;
        RECT  5.185 3.440 6.050 3.940 ;
        RECT  4.925 3.285 5.185 3.940 ;
        RECT  3.395 3.440 4.925 3.940 ;
        RECT  3.135 3.285 3.395 3.940 ;
        RECT  2.595 3.440 3.135 3.940 ;
        RECT  2.335 3.285 2.595 3.940 ;
        RECT  0.795 3.440 2.335 3.940 ;
        RECT  0.535 2.955 0.795 3.940 ;
        RECT  0.000 3.440 0.535 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.875 1.585 11.905 1.845 ;
        RECT  11.715 1.585 11.875 2.755 ;
        RECT  11.175 2.595 11.715 2.755 ;
        RECT  11.455 0.705 11.695 0.965 ;
        RECT  11.435 0.705 11.455 2.205 ;
        RECT  11.295 0.805 11.435 2.205 ;
        RECT  11.265 1.125 11.295 1.385 ;
        RECT  11.195 2.045 11.295 2.205 ;
        RECT  11.015 2.595 11.175 3.065 ;
        RECT  11.085 1.605 11.115 1.865 ;
        RECT  10.925 0.585 11.085 1.865 ;
        RECT  10.915 2.605 11.015 3.065 ;
        RECT  10.205 0.585 10.925 0.745 ;
        RECT  10.745 2.605 10.915 2.765 ;
        RECT  10.585 0.925 10.745 2.765 ;
        RECT  9.865 0.925 10.585 1.085 ;
        RECT  8.185 2.605 10.585 2.765 ;
        RECT  10.245 1.365 10.405 2.425 ;
        RECT  9.325 1.365 10.245 1.525 ;
        RECT  7.935 2.265 10.245 2.425 ;
        RECT  10.045 0.430 10.205 0.745 ;
        RECT  9.865 0.430 10.045 0.650 ;
        RECT  9.285 0.490 9.865 0.650 ;
        RECT  9.605 0.835 9.865 1.085 ;
        RECT  8.735 0.925 9.605 1.085 ;
        RECT  9.065 1.265 9.325 1.525 ;
        RECT  9.125 0.490 9.285 0.745 ;
        RECT  6.935 0.585 9.125 0.745 ;
        RECT  8.395 1.365 9.065 1.525 ;
        RECT  8.575 0.925 8.735 1.185 ;
        RECT  8.235 0.930 8.395 1.525 ;
        RECT  7.920 2.985 8.275 3.145 ;
        RECT  7.195 0.930 8.235 1.090 ;
        RECT  7.885 2.265 7.935 2.525 ;
        RECT  7.760 2.945 7.920 3.145 ;
        RECT  7.675 2.165 7.885 2.525 ;
        RECT  5.770 2.945 7.760 3.105 ;
        RECT  6.975 2.165 7.675 2.325 ;
        RECT  7.025 1.620 7.285 1.920 ;
        RECT  6.265 1.760 7.025 1.920 ;
        RECT  6.715 2.165 6.975 2.765 ;
        RECT  6.775 0.585 6.935 0.930 ;
        RECT  6.015 0.770 6.775 0.930 ;
        RECT  5.925 2.165 6.715 2.325 ;
        RECT  6.105 1.110 6.265 1.920 ;
        RECT  5.815 1.110 6.105 1.270 ;
        RECT  5.755 0.645 6.015 0.930 ;
        RECT  5.765 1.750 5.925 2.325 ;
        RECT  5.585 1.110 5.815 1.285 ;
        RECT  5.510 2.830 5.770 3.105 ;
        RECT  4.125 0.770 5.755 0.930 ;
        RECT  5.425 1.110 5.585 2.640 ;
        RECT  3.935 2.945 5.510 3.105 ;
        RECT  4.305 1.110 5.425 1.270 ;
        RECT  5.305 2.375 5.425 2.640 ;
        RECT  4.275 2.375 5.305 2.535 ;
        RECT  3.960 1.450 5.245 1.610 ;
        RECT  3.785 0.430 4.365 0.590 ;
        RECT  4.115 2.150 4.275 2.750 ;
        RECT  3.965 0.770 4.125 1.090 ;
        RECT  3.015 0.930 3.965 1.090 ;
        RECT  3.935 1.270 3.960 1.610 ;
        RECT  3.775 1.270 3.935 3.105 ;
        RECT  3.625 0.430 3.785 0.750 ;
        RECT  3.195 1.270 3.775 1.430 ;
        RECT  1.645 2.945 3.775 3.105 ;
        RECT  2.675 0.590 3.625 0.750 ;
        RECT  3.435 1.700 3.595 1.960 ;
        RECT  3.015 1.800 3.435 1.960 ;
        RECT  2.995 0.930 3.015 1.960 ;
        RECT  2.855 0.930 2.995 2.760 ;
        RECT  2.825 1.800 2.855 2.760 ;
        RECT  2.735 2.160 2.825 2.760 ;
        RECT  1.475 2.495 2.735 2.655 ;
        RECT  2.515 0.590 2.675 1.355 ;
        RECT  1.845 1.195 2.515 1.355 ;
        RECT  1.820 2.055 2.045 2.315 ;
        RECT  1.820 0.970 1.845 1.355 ;
        RECT  1.660 0.970 1.820 2.315 ;
        RECT  1.655 0.430 1.705 0.690 ;
        RECT  1.585 0.970 1.660 1.230 ;
        RECT  1.445 0.430 1.655 0.745 ;
        RECT  1.385 2.885 1.645 3.145 ;
        RECT  1.315 1.575 1.475 2.655 ;
        RECT  0.795 0.585 1.445 0.745 ;
        RECT  1.135 2.885 1.385 3.045 ;
        RECT  1.135 0.970 1.335 1.230 ;
        RECT  0.975 0.970 1.135 3.045 ;
        RECT  0.635 0.585 0.795 1.080 ;
        RECT  0.385 0.905 0.635 1.080 ;
        RECT  0.285 0.905 0.385 1.165 ;
        RECT  0.285 2.085 0.385 2.345 ;
        RECT  0.125 0.905 0.285 2.345 ;
    END
END DFFRHQX4

MACRO DFFRHQX2
    CLASS CORE ;
    FOREIGN DFFRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.075 1.635 7.335 1.895 ;
        RECT  6.340 1.635 7.075 1.795 ;
        RECT  6.130 1.635 6.340 2.145 ;
        RECT  6.060 1.635 6.130 1.795 ;
        RECT  5.395 1.985 6.130 2.145 ;
        RECT  5.360 1.985 5.395 2.400 ;
        RECT  5.200 1.890 5.360 2.400 ;
        RECT  5.185 2.110 5.200 2.400 ;
        END
        ANTENNAGATEAREA     0.2314 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.735 0.590 9.995 3.040 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.395 1.490 2.655 1.990 ;
        END
        ANTENNAGATEAREA     0.0780 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.495 0.460 1.995 ;
        END
        ANTENNAGATEAREA     0.2444 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.335 -0.250 10.120 0.250 ;
        RECT  9.075 -0.250 9.335 1.295 ;
        RECT  7.650 -0.250 9.075 0.250 ;
        RECT  7.390 -0.250 7.650 0.405 ;
        RECT  4.975 -0.250 7.390 0.250 ;
        RECT  4.715 -0.250 4.975 0.565 ;
        RECT  3.215 -0.250 4.715 0.250 ;
        RECT  2.955 -0.250 3.215 0.405 ;
        RECT  2.425 -0.250 2.955 0.250 ;
        RECT  2.165 -0.250 2.425 0.405 ;
        RECT  0.935 -0.250 2.165 0.250 ;
        RECT  0.675 -0.250 0.935 0.405 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.455 3.440 10.120 3.940 ;
        RECT  9.195 3.285 9.455 3.940 ;
        RECT  8.105 3.440 9.195 3.940 ;
        RECT  7.845 3.065 8.105 3.940 ;
        RECT  6.215 3.440 7.845 3.940 ;
        RECT  5.955 3.285 6.215 3.940 ;
        RECT  5.160 3.440 5.955 3.940 ;
        RECT  4.900 3.285 5.160 3.940 ;
        RECT  3.455 3.440 4.900 3.940 ;
        RECT  2.515 3.285 3.455 3.940 ;
        RECT  0.795 3.440 2.515 3.940 ;
        RECT  0.535 2.825 0.795 3.940 ;
        RECT  0.000 3.440 0.535 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.315 1.485 9.415 1.745 ;
        RECT  9.155 1.485 9.315 2.775 ;
        RECT  8.855 2.615 9.155 2.775 ;
        RECT  8.815 1.830 8.975 2.215 ;
        RECT  8.595 2.615 8.855 3.115 ;
        RECT  8.705 1.830 8.815 1.990 ;
        RECT  8.545 0.485 8.705 1.990 ;
        RECT  8.435 2.170 8.595 2.430 ;
        RECT  8.025 2.615 8.595 2.775 ;
        RECT  8.365 2.170 8.435 2.330 ;
        RECT  8.205 0.585 8.365 2.330 ;
        RECT  7.000 0.585 8.205 0.745 ;
        RECT  7.865 0.955 8.025 2.775 ;
        RECT  6.380 0.955 7.865 1.115 ;
        RECT  7.145 2.615 7.865 2.775 ;
        RECT  7.525 1.295 7.685 2.375 ;
        RECT  6.010 1.295 7.525 1.455 ;
        RECT  6.685 2.160 7.525 2.320 ;
        RECT  6.985 2.505 7.145 2.775 ;
        RECT  6.840 0.470 7.000 0.745 ;
        RECT  6.835 2.955 6.935 3.215 ;
        RECT  6.660 0.470 6.840 0.630 ;
        RECT  6.675 2.945 6.835 3.215 ;
        RECT  6.520 2.160 6.685 2.760 ;
        RECT  4.760 2.945 6.675 3.105 ;
        RECT  6.400 0.430 6.660 0.630 ;
        RECT  6.425 2.500 6.520 2.760 ;
        RECT  4.935 2.600 6.425 2.760 ;
        RECT  5.355 0.470 6.400 0.630 ;
        RECT  6.220 0.855 6.380 1.115 ;
        RECT  5.850 0.810 6.010 1.455 ;
        RECT  5.630 0.810 5.850 1.070 ;
        RECT  5.510 1.405 5.670 1.670 ;
        RECT  5.450 1.405 5.510 1.565 ;
        RECT  5.290 1.225 5.450 1.565 ;
        RECT  5.195 0.470 5.355 0.905 ;
        RECT  4.200 1.225 5.290 1.385 ;
        RECT  4.410 0.745 5.195 0.905 ;
        RECT  4.775 1.595 4.935 2.760 ;
        RECT  4.630 1.595 4.775 1.855 ;
        RECT  4.500 2.945 4.760 3.125 ;
        RECT  3.680 2.945 4.500 3.105 ;
        RECT  4.200 2.500 4.420 2.760 ;
        RECT  4.150 0.645 4.410 0.905 ;
        RECT  4.160 1.225 4.200 2.760 ;
        RECT  4.040 1.175 4.160 2.760 ;
        RECT  2.415 0.745 4.150 0.905 ;
        RECT  4.000 1.175 4.040 1.435 ;
        RECT  3.820 1.545 3.855 1.805 ;
        RECT  3.660 1.085 3.820 1.805 ;
        RECT  3.520 2.150 3.680 3.105 ;
        RECT  2.995 1.085 3.660 1.245 ;
        RECT  3.480 2.150 3.520 2.310 ;
        RECT  1.765 2.945 3.520 3.105 ;
        RECT  3.335 1.605 3.480 2.310 ;
        RECT  2.600 2.605 3.340 2.765 ;
        RECT  3.320 1.555 3.335 2.310 ;
        RECT  3.175 1.555 3.320 1.815 ;
        RECT  2.995 2.225 3.140 2.385 ;
        RECT  2.835 1.085 2.995 2.385 ;
        RECT  2.595 1.085 2.835 1.245 ;
        RECT  2.440 2.245 2.600 2.765 ;
        RECT  2.200 2.245 2.440 2.405 ;
        RECT  2.255 0.745 2.415 1.145 ;
        RECT  1.825 0.985 2.255 1.145 ;
        RECT  2.100 2.145 2.200 2.405 ;
        RECT  1.940 1.990 2.100 2.405 ;
        RECT  1.475 0.605 2.045 0.765 ;
        RECT  1.825 1.990 1.940 2.150 ;
        RECT  1.665 0.985 1.825 2.150 ;
        RECT  1.665 2.660 1.765 3.105 ;
        RECT  1.335 1.890 1.665 2.150 ;
        RECT  1.605 2.415 1.665 3.105 ;
        RECT  1.505 2.415 1.605 2.920 ;
        RECT  1.140 2.415 1.505 2.575 ;
        RECT  1.315 0.585 1.475 0.765 ;
        RECT  1.140 1.035 1.365 1.295 ;
        RECT  0.800 0.585 1.315 0.745 ;
        RECT  0.980 1.035 1.140 2.575 ;
        RECT  0.640 0.585 0.800 2.335 ;
        RECT  0.125 1.035 0.640 1.295 ;
        RECT  0.385 2.175 0.640 2.335 ;
        RECT  0.125 2.175 0.385 2.435 ;
    END
END DFFRHQX2

MACRO DFFRHQX1
    CLASS CORE ;
    FOREIGN DFFRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.895 1.605 7.055 1.955 ;
        RECT  5.395 1.795 6.895 1.955 ;
        RECT  5.185 1.700 5.395 1.990 ;
        RECT  5.035 1.795 5.185 1.955 ;
        END
        ANTENNAGATEAREA     0.1430 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.375 0.970 9.535 2.580 ;
        RECT  9.275 0.970 9.375 1.230 ;
        RECT  9.275 1.980 9.375 2.580 ;
        END
        ANTENNADIFFAREA     0.3944 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.290 1.945 1.615 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.495 0.395 1.995 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.995 -0.250 9.660 0.250 ;
        RECT  8.735 -0.250 8.995 0.840 ;
        RECT  7.625 -0.250 8.735 0.250 ;
        RECT  7.365 -0.250 7.625 0.405 ;
        RECT  4.975 -0.250 7.365 0.250 ;
        RECT  4.715 -0.250 4.975 0.405 ;
        RECT  3.365 -0.250 4.715 0.250 ;
        RECT  3.105 -0.250 3.365 0.405 ;
        RECT  1.320 -0.250 3.105 0.250 ;
        RECT  0.720 -0.250 1.320 0.405 ;
        RECT  0.000 -0.250 0.720 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.985 3.440 9.660 3.940 ;
        RECT  8.725 3.285 8.985 3.940 ;
        RECT  7.420 3.440 8.725 3.940 ;
        RECT  7.160 3.065 7.420 3.940 ;
        RECT  5.845 3.440 7.160 3.940 ;
        RECT  5.585 3.285 5.845 3.940 ;
        RECT  5.080 3.440 5.585 3.940 ;
        RECT  4.820 3.285 5.080 3.940 ;
        RECT  3.410 3.440 4.820 3.940 ;
        RECT  3.150 3.285 3.410 3.940 ;
        RECT  2.350 3.440 3.150 3.940 ;
        RECT  2.090 3.285 2.350 3.940 ;
        RECT  0.820 3.440 2.090 3.940 ;
        RECT  0.560 2.755 0.820 3.940 ;
        RECT  0.000 3.440 0.560 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.875 1.485 9.195 1.745 ;
        RECT  8.715 1.485 8.875 2.825 ;
        RECT  8.595 1.485 8.715 1.745 ;
        RECT  8.310 2.665 8.715 2.825 ;
        RECT  8.415 1.980 8.470 2.240 ;
        RECT  8.415 1.035 8.440 1.320 ;
        RECT  8.255 0.485 8.415 2.240 ;
        RECT  8.050 2.665 8.310 3.000 ;
        RECT  7.915 0.585 8.075 2.485 ;
        RECT  7.735 2.665 8.050 2.825 ;
        RECT  7.050 0.585 7.915 0.745 ;
        RECT  7.575 0.925 7.735 2.825 ;
        RECT  6.335 0.925 7.575 1.085 ;
        RECT  6.925 2.665 7.575 2.825 ;
        RECT  7.235 1.265 7.395 2.295 ;
        RECT  5.995 1.265 7.235 1.425 ;
        RECT  6.415 2.135 7.235 2.295 ;
        RECT  6.890 0.470 7.050 0.745 ;
        RECT  6.665 2.500 6.925 2.825 ;
        RECT  6.185 0.470 6.890 0.630 ;
        RECT  6.370 2.945 6.530 3.215 ;
        RECT  6.155 2.135 6.415 2.765 ;
        RECT  3.800 2.945 6.370 3.105 ;
        RECT  6.175 0.810 6.335 1.085 ;
        RECT  5.925 0.445 6.185 0.630 ;
        RECT  5.440 2.605 6.155 2.765 ;
        RECT  5.835 0.910 5.995 1.425 ;
        RECT  5.340 0.470 5.925 0.630 ;
        RECT  5.575 0.810 5.835 1.070 ;
        RECT  5.455 1.265 5.615 1.525 ;
        RECT  4.140 1.285 5.455 1.445 ;
        RECT  5.180 2.175 5.440 2.765 ;
        RECT  5.180 0.470 5.340 1.105 ;
        RECT  4.435 0.945 5.180 1.105 ;
        RECT  4.730 2.605 5.180 2.765 ;
        RECT  4.730 1.625 4.745 1.785 ;
        RECT  4.570 1.625 4.730 2.765 ;
        RECT  4.485 1.625 4.570 1.785 ;
        RECT  4.175 0.650 4.435 1.105 ;
        RECT  3.680 0.945 4.175 1.105 ;
        RECT  3.980 1.285 4.140 2.690 ;
        RECT  3.970 1.285 3.980 1.445 ;
        RECT  3.745 0.475 3.905 0.765 ;
        RECT  3.640 1.625 3.800 3.105 ;
        RECT  3.315 0.605 3.745 0.765 ;
        RECT  3.520 0.945 3.680 1.375 ;
        RECT  3.465 1.625 3.640 1.785 ;
        RECT  1.160 2.945 3.640 3.105 ;
        RECT  2.735 1.215 3.520 1.375 ;
        RECT  3.205 1.555 3.465 1.785 ;
        RECT  3.300 2.035 3.460 2.295 ;
        RECT  3.155 0.605 3.315 1.035 ;
        RECT  2.735 2.135 3.300 2.295 ;
        RECT  2.300 0.875 3.155 1.035 ;
        RECT  1.660 0.535 2.975 0.695 ;
        RECT  2.735 2.505 2.860 2.765 ;
        RECT  2.575 1.215 2.735 2.765 ;
        RECT  1.515 2.605 2.575 2.765 ;
        RECT  2.140 0.875 2.300 2.425 ;
        RECT  1.840 0.875 2.140 1.035 ;
        RECT  1.500 0.535 1.660 0.745 ;
        RECT  1.355 1.815 1.515 2.765 ;
        RECT  0.735 0.585 1.500 0.745 ;
        RECT  1.075 0.950 1.410 1.110 ;
        RECT  1.300 1.815 1.355 2.075 ;
        RECT  1.075 2.260 1.160 3.105 ;
        RECT  1.000 0.950 1.075 3.105 ;
        RECT  0.915 0.950 1.000 2.420 ;
        RECT  0.575 0.585 0.735 2.345 ;
        RECT  0.140 1.035 0.575 1.295 ;
        RECT  0.400 2.185 0.575 2.345 ;
        RECT  0.140 2.185 0.400 2.445 ;
    END
END DFFRHQX1

MACRO DFFHQX8
    CLASS CORE ;
    FOREIGN DFFHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.340 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.650 1.515 12.755 1.765 ;
        RECT  12.390 0.595 12.650 3.055 ;
        RECT  11.630 1.700 12.390 2.400 ;
        RECT  11.370 0.595 11.630 3.055 ;
        END
        ANTENNADIFFAREA     1.6264 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 1.290 2.635 1.580 ;
        RECT  2.125 1.290 2.485 1.695 ;
        END
        ANTENNAGATEAREA     0.1443 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 1.455 0.825 2.015 ;
        END
        ANTENNAGATEAREA     0.3731 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.160 -0.250 13.340 0.250 ;
        RECT  12.900 -0.250 13.160 1.095 ;
        RECT  12.140 -0.250 12.900 0.250 ;
        RECT  11.880 -0.250 12.140 1.095 ;
        RECT  11.120 -0.250 11.880 0.250 ;
        RECT  10.860 -0.250 11.120 0.755 ;
        RECT  10.150 -0.250 10.860 0.250 ;
        RECT  9.890 -0.250 10.150 0.950 ;
        RECT  7.430 -0.250 9.890 0.250 ;
        RECT  7.170 -0.250 7.430 0.405 ;
        RECT  6.490 -0.250 7.170 0.250 ;
        RECT  6.230 -0.250 6.490 0.405 ;
        RECT  5.375 -0.250 6.230 0.250 ;
        RECT  5.115 -0.250 5.375 0.405 ;
        RECT  3.785 -0.250 5.115 0.250 ;
        RECT  3.625 -0.250 3.785 1.070 ;
        RECT  2.455 -0.250 3.625 0.250 ;
        RECT  3.435 0.810 3.625 1.070 ;
        RECT  2.295 -0.250 2.455 0.735 ;
        RECT  0.785 -0.250 2.295 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.160 3.440 13.340 3.940 ;
        RECT  12.900 2.275 13.160 3.940 ;
        RECT  12.140 3.440 12.900 3.940 ;
        RECT  11.880 2.615 12.140 3.940 ;
        RECT  11.120 3.440 11.880 3.940 ;
        RECT  10.520 2.955 11.120 3.940 ;
        RECT  7.470 3.440 10.520 3.940 ;
        RECT  7.210 3.285 7.470 3.940 ;
        RECT  6.390 3.440 7.210 3.940 ;
        RECT  6.130 3.285 6.390 3.940 ;
        RECT  4.755 3.440 6.130 3.940 ;
        RECT  4.495 3.285 4.755 3.940 ;
        RECT  3.395 3.440 4.495 3.940 ;
        RECT  3.135 3.285 3.395 3.940 ;
        RECT  2.445 3.440 3.135 3.940 ;
        RECT  2.185 3.285 2.445 3.940 ;
        RECT  0.825 3.440 2.185 3.940 ;
        RECT  0.565 2.955 0.825 3.940 ;
        RECT  0.000 3.440 0.565 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.050 1.510 11.100 1.770 ;
        RECT  10.890 1.510 11.050 2.730 ;
        RECT  10.840 1.510 10.890 1.770 ;
        RECT  9.740 2.570 10.890 2.730 ;
        RECT  10.610 1.035 10.660 1.295 ;
        RECT  10.610 2.040 10.660 2.300 ;
        RECT  10.450 1.035 10.610 2.300 ;
        RECT  10.400 1.035 10.450 1.295 ;
        RECT  10.030 1.500 10.450 1.760 ;
        RECT  10.400 2.040 10.450 2.300 ;
        RECT  9.720 2.065 9.980 2.325 ;
        RECT  9.300 2.505 9.740 2.765 ;
        RECT  9.700 2.065 9.720 2.225 ;
        RECT  9.540 0.570 9.700 2.225 ;
        RECT  9.400 2.945 9.660 3.220 ;
        RECT  9.450 0.570 9.540 0.730 ;
        RECT  9.190 0.470 9.450 0.730 ;
        RECT  5.980 2.945 9.400 3.105 ;
        RECT  9.200 1.200 9.360 1.530 ;
        RECT  9.140 2.165 9.300 2.765 ;
        RECT  8.450 1.200 9.200 1.360 ;
        RECT  7.770 0.470 9.190 0.630 ;
        RECT  8.450 2.165 9.140 2.325 ;
        RECT  8.110 0.810 9.010 0.970 ;
        RECT  8.630 2.505 8.890 2.765 ;
        RECT  7.870 2.605 8.630 2.765 ;
        RECT  8.380 1.150 8.450 2.325 ;
        RECT  8.290 1.150 8.380 2.425 ;
        RECT  8.120 2.165 8.290 2.425 ;
        RECT  7.950 0.810 8.110 1.085 ;
        RECT  7.940 0.925 7.950 1.085 ;
        RECT  7.680 0.925 7.940 1.185 ;
        RECT  7.610 2.505 7.870 2.765 ;
        RECT  7.610 0.470 7.770 0.745 ;
        RECT  7.100 0.925 7.680 1.085 ;
        RECT  4.815 0.585 7.610 0.745 ;
        RECT  6.930 2.605 7.610 2.765 ;
        RECT  6.940 0.925 7.100 2.170 ;
        RECT  6.770 0.925 6.940 1.185 ;
        RECT  6.930 2.010 6.940 2.170 ;
        RECT  6.670 2.010 6.930 2.765 ;
        RECT  6.590 1.515 6.760 1.775 ;
        RECT  6.250 2.010 6.670 2.170 ;
        RECT  6.430 0.955 6.590 1.775 ;
        RECT  5.700 0.955 6.430 1.115 ;
        RECT  6.090 1.535 6.250 2.170 ;
        RECT  5.990 1.535 6.090 1.795 ;
        RECT  5.720 2.845 5.980 3.105 ;
        RECT  3.335 2.945 5.720 3.105 ;
        RECT  5.510 0.925 5.700 1.115 ;
        RECT  5.510 2.405 5.610 2.665 ;
        RECT  5.350 0.925 5.510 2.665 ;
        RECT  4.475 0.925 5.350 1.085 ;
        RECT  3.905 2.405 5.350 2.565 ;
        RECT  4.655 0.470 4.815 0.745 ;
        RECT  4.405 1.905 4.665 2.165 ;
        RECT  4.135 0.470 4.655 0.630 ;
        RECT  4.315 0.810 4.475 1.085 ;
        RECT  4.135 1.905 4.405 2.065 ;
        RECT  3.975 0.470 4.135 2.065 ;
        RECT  3.135 1.250 3.975 1.445 ;
        RECT  3.645 2.405 3.905 2.760 ;
        RECT  3.385 1.625 3.645 1.885 ;
        RECT  2.795 0.470 3.445 0.630 ;
        RECT  3.335 1.725 3.385 1.885 ;
        RECT  3.175 1.725 3.335 3.105 ;
        RECT  1.645 2.945 3.175 3.105 ;
        RECT  2.995 0.810 3.135 1.445 ;
        RECT  2.975 0.810 2.995 2.765 ;
        RECT  2.835 1.285 2.975 2.765 ;
        RECT  2.735 2.165 2.835 2.765 ;
        RECT  2.635 0.470 2.795 1.085 ;
        RECT  1.605 2.605 2.735 2.765 ;
        RECT  1.965 0.925 2.635 1.085 ;
        RECT  1.945 2.165 2.045 2.425 ;
        RECT  1.945 0.925 1.965 1.185 ;
        RECT  1.785 0.925 1.945 2.425 ;
        RECT  1.705 0.925 1.785 1.185 ;
        RECT  1.445 0.485 1.705 0.745 ;
        RECT  1.385 2.945 1.645 3.205 ;
        RECT  1.445 1.585 1.605 2.765 ;
        RECT  0.385 0.585 1.445 0.745 ;
        RECT  1.345 1.585 1.445 1.845 ;
        RECT  1.165 2.945 1.385 3.105 ;
        RECT  1.165 0.970 1.335 1.230 ;
        RECT  1.005 0.970 1.165 3.105 ;
        RECT  0.365 0.585 0.385 1.165 ;
        RECT  0.365 2.225 0.385 2.485 ;
        RECT  0.225 0.585 0.365 2.485 ;
        RECT  0.205 0.905 0.225 2.485 ;
        RECT  0.125 0.905 0.205 1.165 ;
        RECT  0.125 2.225 0.205 2.485 ;
    END
END DFFHQX8

MACRO DFFHQX4
    CLASS CORE ;
    FOREIGN DFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.420 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.740 1.515 11.835 2.585 ;
        RECT  11.480 0.600 11.740 3.050 ;
        END
        ANTENNADIFFAREA     0.8132 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.525 2.635 1.990 ;
        RECT  2.225 1.525 2.425 1.820 ;
        END
        ANTENNAGATEAREA     0.1443 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.525 1.290 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.3731 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.250 -0.250 12.420 0.250 ;
        RECT  11.990 -0.250 12.250 1.095 ;
        RECT  11.230 -0.250 11.990 0.250 ;
        RECT  10.970 -0.250 11.230 0.755 ;
        RECT  10.245 -0.250 10.970 0.250 ;
        RECT  9.985 -0.250 10.245 0.950 ;
        RECT  7.470 -0.250 9.985 0.250 ;
        RECT  7.210 -0.250 7.470 0.405 ;
        RECT  6.530 -0.250 7.210 0.250 ;
        RECT  6.270 -0.250 6.530 0.405 ;
        RECT  5.425 -0.250 6.270 0.250 ;
        RECT  5.165 -0.250 5.425 0.405 ;
        RECT  3.785 -0.250 5.165 0.250 ;
        RECT  3.625 -0.250 3.785 1.070 ;
        RECT  2.455 -0.250 3.625 0.250 ;
        RECT  3.435 0.810 3.625 1.070 ;
        RECT  2.295 -0.250 2.455 0.965 ;
        RECT  0.875 -0.250 2.295 0.250 ;
        RECT  0.615 -0.250 0.875 0.405 ;
        RECT  0.000 -0.250 0.615 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.275 3.440 12.420 3.940 ;
        RECT  12.015 2.275 12.275 3.940 ;
        RECT  11.230 3.440 12.015 3.940 ;
        RECT  10.630 2.955 11.230 3.940 ;
        RECT  7.525 3.440 10.630 3.940 ;
        RECT  7.265 3.285 7.525 3.940 ;
        RECT  6.435 3.440 7.265 3.940 ;
        RECT  6.175 3.285 6.435 3.940 ;
        RECT  4.845 3.440 6.175 3.940 ;
        RECT  4.585 3.285 4.845 3.940 ;
        RECT  3.485 3.440 4.585 3.940 ;
        RECT  3.225 3.285 3.485 3.940 ;
        RECT  2.685 3.440 3.225 3.940 ;
        RECT  2.425 3.285 2.685 3.940 ;
        RECT  0.915 3.440 2.425 3.940 ;
        RECT  0.655 2.880 0.915 3.940 ;
        RECT  0.000 3.440 0.655 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.115 1.510 11.215 1.770 ;
        RECT  10.955 1.510 11.115 2.670 ;
        RECT  9.795 2.510 10.955 2.670 ;
        RECT  10.705 1.035 10.755 1.295 ;
        RECT  10.705 2.040 10.745 2.300 ;
        RECT  10.545 1.035 10.705 2.300 ;
        RECT  10.495 1.035 10.545 1.295 ;
        RECT  10.230 1.540 10.545 1.700 ;
        RECT  10.485 2.040 10.545 2.300 ;
        RECT  9.970 1.490 10.230 1.750 ;
        RECT  9.790 1.970 10.025 2.230 ;
        RECT  9.355 2.410 9.795 2.670 ;
        RECT  9.630 0.570 9.790 2.230 ;
        RECT  9.455 2.945 9.715 3.260 ;
        RECT  9.540 0.570 9.630 0.730 ;
        RECT  9.280 0.470 9.540 0.730 ;
        RECT  6.065 2.945 9.455 3.105 ;
        RECT  9.290 1.150 9.450 1.530 ;
        RECT  9.195 2.165 9.355 2.670 ;
        RECT  8.490 1.150 9.290 1.310 ;
        RECT  7.810 0.470 9.280 0.630 ;
        RECT  8.490 2.165 9.195 2.325 ;
        RECT  8.150 0.810 9.100 0.970 ;
        RECT  8.685 2.505 8.945 2.765 ;
        RECT  7.925 2.605 8.685 2.765 ;
        RECT  8.435 1.150 8.490 2.325 ;
        RECT  8.330 1.150 8.435 2.425 ;
        RECT  8.175 2.165 8.330 2.425 ;
        RECT  7.990 0.810 8.150 1.085 ;
        RECT  7.980 0.925 7.990 1.085 ;
        RECT  7.720 0.925 7.980 1.185 ;
        RECT  7.665 2.360 7.925 2.765 ;
        RECT  7.650 0.470 7.810 0.745 ;
        RECT  7.495 0.925 7.720 1.085 ;
        RECT  6.985 2.605 7.665 2.765 ;
        RECT  5.985 0.585 7.650 0.745 ;
        RECT  7.335 0.925 7.495 2.170 ;
        RECT  7.070 0.925 7.335 1.135 ;
        RECT  6.985 2.010 7.335 2.170 ;
        RECT  6.630 1.515 7.155 1.775 ;
        RECT  6.810 0.925 7.070 1.185 ;
        RECT  6.725 2.010 6.985 2.765 ;
        RECT  6.290 2.010 6.725 2.170 ;
        RECT  6.470 1.025 6.630 1.775 ;
        RECT  5.785 1.025 6.470 1.185 ;
        RECT  6.130 1.535 6.290 2.170 ;
        RECT  6.030 1.535 6.130 1.795 ;
        RECT  5.805 2.845 6.065 3.105 ;
        RECT  5.725 0.435 5.985 0.745 ;
        RECT  3.555 2.945 5.805 3.105 ;
        RECT  5.495 0.925 5.785 1.185 ;
        RECT  4.985 0.585 5.725 0.745 ;
        RECT  5.495 2.305 5.695 2.565 ;
        RECT  5.335 0.925 5.495 2.695 ;
        RECT  4.565 0.925 5.335 1.085 ;
        RECT  3.995 2.535 5.335 2.695 ;
        RECT  4.825 0.565 4.985 0.745 ;
        RECT  4.125 0.565 4.825 0.725 ;
        RECT  4.615 1.925 4.665 2.185 ;
        RECT  4.405 1.905 4.615 2.185 ;
        RECT  4.305 0.905 4.565 1.165 ;
        RECT  4.125 1.905 4.405 2.065 ;
        RECT  3.965 0.565 4.125 2.065 ;
        RECT  3.735 2.485 3.995 2.745 ;
        RECT  3.215 1.250 3.965 1.410 ;
        RECT  3.555 1.590 3.785 1.850 ;
        RECT  3.395 1.590 3.555 3.105 ;
        RECT  2.795 0.470 3.445 0.630 ;
        RECT  1.735 2.945 3.395 3.105 ;
        RECT  3.135 1.250 3.215 2.325 ;
        RECT  3.085 1.030 3.135 2.325 ;
        RECT  3.055 1.030 3.085 2.765 ;
        RECT  2.975 1.030 3.055 1.410 ;
        RECT  2.825 2.165 3.055 2.765 ;
        RECT  1.635 2.500 2.825 2.660 ;
        RECT  2.635 0.470 2.795 1.305 ;
        RECT  2.035 1.145 2.635 1.305 ;
        RECT  2.035 2.060 2.135 2.320 ;
        RECT  1.965 1.145 2.035 2.320 ;
        RECT  1.875 0.960 1.965 2.320 ;
        RECT  1.705 0.960 1.875 1.305 ;
        RECT  1.565 0.520 1.825 0.780 ;
        RECT  1.475 2.845 1.735 3.105 ;
        RECT  1.475 1.585 1.635 2.660 ;
        RECT  0.475 0.620 1.565 0.780 ;
        RECT  1.315 1.585 1.475 1.845 ;
        RECT  1.255 2.845 1.475 3.005 ;
        RECT  1.165 0.960 1.425 1.295 ;
        RECT  1.135 2.150 1.255 3.005 ;
        RECT  1.135 1.135 1.165 1.295 ;
        RECT  1.095 1.135 1.135 3.005 ;
        RECT  0.975 1.135 1.095 2.310 ;
        RECT  0.340 0.620 0.475 1.035 ;
        RECT  0.340 2.225 0.475 2.485 ;
        RECT  0.180 0.620 0.340 2.485 ;
    END
END DFFHQX4

MACRO DFFHQX2
    CLASS CORE ;
    FOREIGN DFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.525 0.695 9.535 2.995 ;
        RECT  9.325 0.590 9.525 3.055 ;
        RECT  9.265 0.590 9.325 1.290 ;
        RECT  9.315 1.765 9.325 3.055 ;
        RECT  9.265 2.115 9.315 3.055 ;
        END
        ANTENNADIFFAREA     0.7276 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.265 1.410 2.365 1.670 ;
        RECT  1.990 1.410 2.265 1.990 ;
        RECT  1.965 1.700 1.990 1.990 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.475 0.920 1.990 ;
        END
        ANTENNAGATEAREA     0.2353 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.015 -0.250 9.660 0.250 ;
        RECT  8.755 -0.250 9.015 1.095 ;
        RECT  7.725 -0.250 8.755 0.250 ;
        RECT  7.465 -0.250 7.725 1.045 ;
        RECT  5.675 -0.250 7.465 0.250 ;
        RECT  5.415 -0.250 5.675 0.405 ;
        RECT  4.535 -0.250 5.415 0.250 ;
        RECT  4.275 -0.250 4.535 0.405 ;
        RECT  2.415 -0.250 4.275 0.250 ;
        RECT  2.255 -0.250 2.415 0.625 ;
        RECT  0.815 -0.250 2.255 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.015 3.440 9.660 3.940 ;
        RECT  8.415 2.795 9.015 3.940 ;
        RECT  6.055 3.440 8.415 3.940 ;
        RECT  5.795 3.285 6.055 3.940 ;
        RECT  5.105 3.440 5.795 3.940 ;
        RECT  4.845 3.285 5.105 3.940 ;
        RECT  3.655 3.440 4.845 3.940 ;
        RECT  3.395 3.285 3.655 3.940 ;
        RECT  2.595 3.440 3.395 3.940 ;
        RECT  2.335 3.285 2.595 3.940 ;
        RECT  0.855 3.440 2.335 3.940 ;
        RECT  0.595 2.695 0.855 3.940 ;
        RECT  0.000 3.440 0.595 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.905 1.510 8.965 1.770 ;
        RECT  8.745 1.510 8.905 2.575 ;
        RECT  8.705 1.510 8.745 1.770 ;
        RECT  7.585 2.415 8.745 2.575 ;
        RECT  8.420 1.955 8.525 2.215 ;
        RECT  8.420 1.035 8.425 1.295 ;
        RECT  8.260 1.035 8.420 2.215 ;
        RECT  8.165 1.035 8.260 1.675 ;
        RECT  8.065 1.415 8.165 1.675 ;
        RECT  7.635 1.225 7.795 2.045 ;
        RECT  7.080 1.225 7.635 1.385 ;
        RECT  7.415 2.225 7.585 2.575 ;
        RECT  7.255 1.615 7.415 2.665 ;
        RECT  6.740 1.615 7.255 1.775 ;
        RECT  6.565 2.505 7.255 2.665 ;
        RECT  7.000 0.585 7.080 1.385 ;
        RECT  6.815 1.955 7.075 2.325 ;
        RECT  6.920 0.430 7.000 1.385 ;
        RECT  6.740 0.430 6.920 0.745 ;
        RECT  6.855 2.845 6.905 3.005 ;
        RECT  6.645 2.845 6.855 3.105 ;
        RECT  6.265 1.955 6.815 2.115 ;
        RECT  5.135 0.585 6.740 0.745 ;
        RECT  6.580 0.925 6.740 1.775 ;
        RECT  4.735 2.945 6.645 3.105 ;
        RECT  6.480 0.925 6.580 1.185 ;
        RECT  6.305 2.295 6.565 2.665 ;
        RECT  6.105 0.925 6.265 2.115 ;
        RECT  5.970 0.925 6.105 1.185 ;
        RECT  5.655 1.955 6.105 2.115 ;
        RECT  5.665 1.515 5.925 1.775 ;
        RECT  5.385 1.515 5.665 1.675 ;
        RECT  5.495 1.955 5.655 2.765 ;
        RECT  5.395 2.165 5.495 2.765 ;
        RECT  5.045 2.165 5.395 2.325 ;
        RECT  5.225 1.150 5.385 1.675 ;
        RECT  4.935 1.150 5.225 1.310 ;
        RECT  4.875 0.485 5.135 0.745 ;
        RECT  4.885 1.515 5.045 2.325 ;
        RECT  4.675 0.925 4.935 1.310 ;
        RECT  4.785 1.515 4.885 1.675 ;
        RECT  4.185 0.585 4.875 0.745 ;
        RECT  4.525 2.805 4.735 3.105 ;
        RECT  4.115 1.150 4.675 1.310 ;
        RECT  4.475 2.805 4.525 3.080 ;
        RECT  1.835 2.920 4.475 3.080 ;
        RECT  4.115 2.025 4.365 2.625 ;
        RECT  4.025 0.585 4.185 0.970 ;
        RECT  4.105 1.150 4.115 2.625 ;
        RECT  3.955 1.150 4.105 2.315 ;
        RECT  3.095 0.810 4.025 0.970 ;
        RECT  3.395 1.150 3.955 1.310 ;
        RECT  3.095 1.645 3.545 1.905 ;
        RECT  2.755 0.470 3.360 0.630 ;
        RECT  3.095 2.140 3.145 2.740 ;
        RECT  2.935 0.810 3.095 2.740 ;
        RECT  2.885 2.140 2.935 2.740 ;
        RECT  1.600 2.530 2.885 2.690 ;
        RECT  2.705 0.470 2.755 1.180 ;
        RECT  2.595 0.470 2.705 2.350 ;
        RECT  2.545 1.020 2.595 2.350 ;
        RECT  2.035 1.020 2.545 1.180 ;
        RECT  1.935 2.190 2.545 2.350 ;
        RECT  1.775 0.970 2.035 1.230 ;
        RECT  1.665 0.470 1.925 0.790 ;
        RECT  1.575 2.870 1.835 3.130 ;
        RECT  0.405 0.630 1.665 0.790 ;
        RECT  1.440 1.695 1.600 2.690 ;
        RECT  1.260 2.920 1.575 3.080 ;
        RECT  1.365 1.035 1.415 1.295 ;
        RECT  1.260 1.030 1.365 1.295 ;
        RECT  1.100 1.030 1.260 3.080 ;
        RECT  0.355 0.630 0.405 1.295 ;
        RECT  0.355 2.075 0.405 2.335 ;
        RECT  0.245 0.630 0.355 2.335 ;
        RECT  0.195 1.035 0.245 2.335 ;
        RECT  0.145 1.035 0.195 1.295 ;
        RECT  0.145 2.075 0.195 2.335 ;
    END
END DFFHQX2

MACRO DFFHQX1
    CLASS CORE ;
    FOREIGN DFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.525 1.105 9.535 2.175 ;
        RECT  9.325 0.975 9.525 2.555 ;
        RECT  9.265 0.975 9.325 1.235 ;
        RECT  9.265 1.955 9.325 2.555 ;
        END
        ANTENNADIFFAREA     0.3944 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.175 1.580 ;
        RECT  1.640 1.290 1.965 1.550 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.695 0.395 1.955 ;
        RECT  0.120 1.520 0.345 2.130 ;
        END
        ANTENNAGATEAREA     0.1456 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.015 -0.250 9.660 0.250 ;
        RECT  8.755 -0.250 9.015 1.235 ;
        RECT  7.825 -0.250 8.755 0.250 ;
        RECT  7.565 -0.250 7.825 1.045 ;
        RECT  5.885 -0.250 7.565 0.250 ;
        RECT  5.625 -0.250 5.885 0.405 ;
        RECT  4.635 -0.250 5.625 0.250 ;
        RECT  4.375 -0.250 4.635 0.405 ;
        RECT  2.635 -0.250 4.375 0.250 ;
        RECT  2.475 -0.250 2.635 0.745 ;
        RECT  1.305 -0.250 2.475 0.250 ;
        RECT  0.705 -0.250 1.305 0.405 ;
        RECT  0.000 -0.250 0.705 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.965 3.440 9.660 3.940 ;
        RECT  8.365 2.895 8.965 3.940 ;
        RECT  6.125 3.440 8.365 3.940 ;
        RECT  5.065 3.285 6.125 3.940 ;
        RECT  3.565 3.440 5.065 3.940 ;
        RECT  3.305 3.285 3.565 3.940 ;
        RECT  2.680 3.440 3.305 3.940 ;
        RECT  2.420 3.285 2.680 3.940 ;
        RECT  0.750 3.440 2.420 3.940 ;
        RECT  0.490 3.285 0.750 3.940 ;
        RECT  0.000 3.440 0.490 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.910 1.510 9.145 1.770 ;
        RECT  8.750 1.510 8.910 2.555 ;
        RECT  8.545 1.510 8.750 1.770 ;
        RECT  7.655 2.395 8.750 2.555 ;
        RECT  8.365 1.955 8.535 2.215 ;
        RECT  8.365 1.035 8.425 1.295 ;
        RECT  8.205 1.035 8.365 2.215 ;
        RECT  8.165 1.035 8.205 1.665 ;
        RECT  8.065 1.405 8.165 1.665 ;
        RECT  7.635 1.225 7.795 2.015 ;
        RECT  7.435 2.245 7.655 2.555 ;
        RECT  7.285 1.225 7.635 1.385 ;
        RECT  7.275 1.565 7.435 2.725 ;
        RECT  7.125 0.635 7.285 1.385 ;
        RECT  6.945 1.565 7.275 1.725 ;
        RECT  6.635 2.565 7.275 2.725 ;
        RECT  6.780 0.635 7.125 0.795 ;
        RECT  6.935 1.905 7.095 2.385 ;
        RECT  6.715 2.905 6.975 3.165 ;
        RECT  6.785 1.025 6.945 1.725 ;
        RECT  6.475 1.905 6.935 2.065 ;
        RECT  6.685 1.025 6.785 1.285 ;
        RECT  6.520 0.585 6.780 0.845 ;
        RECT  4.635 2.905 6.715 3.065 ;
        RECT  6.475 2.245 6.635 2.725 ;
        RECT  5.345 0.635 6.520 0.795 ;
        RECT  6.315 1.025 6.475 2.065 ;
        RECT  6.375 2.245 6.475 2.505 ;
        RECT  6.175 1.025 6.315 1.285 ;
        RECT  5.725 1.905 6.315 2.065 ;
        RECT  5.875 1.465 6.135 1.725 ;
        RECT  5.695 1.465 5.875 1.625 ;
        RECT  5.465 1.905 5.725 2.480 ;
        RECT  5.535 1.150 5.695 1.625 ;
        RECT  5.145 1.150 5.535 1.310 ;
        RECT  5.170 1.905 5.465 2.065 ;
        RECT  5.085 0.595 5.345 0.855 ;
        RECT  5.010 1.515 5.170 2.065 ;
        RECT  4.885 1.035 5.145 1.310 ;
        RECT  4.435 0.635 5.085 0.795 ;
        RECT  4.775 1.515 5.010 1.675 ;
        RECT  4.115 1.150 4.885 1.310 ;
        RECT  4.375 2.785 4.635 3.105 ;
        RECT  4.275 0.635 4.435 0.970 ;
        RECT  4.175 2.155 4.435 2.540 ;
        RECT  1.260 2.945 4.375 3.105 ;
        RECT  3.435 0.810 4.275 0.970 ;
        RECT  4.115 2.155 4.175 2.315 ;
        RECT  3.955 1.150 4.115 2.315 ;
        RECT  2.975 0.470 4.095 0.630 ;
        RECT  3.665 1.150 3.955 1.310 ;
        RECT  3.435 1.785 3.775 2.045 ;
        RECT  3.275 0.810 3.435 2.330 ;
        RECT  3.155 1.035 3.275 1.295 ;
        RECT  3.205 2.170 3.275 2.330 ;
        RECT  3.045 2.170 3.205 2.765 ;
        RECT  2.945 2.345 3.045 2.765 ;
        RECT  2.815 0.470 2.975 1.090 ;
        RECT  1.700 2.605 2.945 2.765 ;
        RECT  2.730 0.930 2.815 1.090 ;
        RECT  2.570 0.930 2.730 2.325 ;
        RECT  1.915 0.930 2.570 1.090 ;
        RECT  2.170 2.165 2.570 2.325 ;
        RECT  2.030 0.450 2.290 0.730 ;
        RECT  1.910 2.165 2.170 2.425 ;
        RECT  1.720 0.570 2.030 0.730 ;
        RECT  1.560 0.570 1.720 1.005 ;
        RECT  1.440 2.345 1.700 2.765 ;
        RECT  0.770 0.845 1.560 1.005 ;
        RECT  1.260 1.185 1.405 1.445 ;
        RECT  1.100 1.185 1.260 3.105 ;
        RECT  0.610 0.845 0.770 2.815 ;
        RECT  0.125 1.035 0.610 1.295 ;
        RECT  0.385 2.655 0.610 2.815 ;
        RECT  0.125 2.655 0.385 2.915 ;
    END
END DFFHQX1

MACRO SEDFFTRX4
    CLASS CORE ;
    FOREIGN SEDFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.320 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.775 1.010 1.935 1.495 ;
        RECT  1.715 1.010 1.775 1.170 ;
        RECT  1.505 0.880 1.715 1.170 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.910 1.700 1.255 2.080 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 0.635 0.335 1.170 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.480 1.085 17.605 1.340 ;
        RECT  17.220 1.085 17.480 2.410 ;
        RECT  17.145 1.290 17.220 2.175 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.560 0.595 18.750 2.335 ;
        RECT  18.525 0.595 18.560 2.400 ;
        RECT  18.425 0.595 18.525 1.195 ;
        RECT  18.500 2.025 18.525 2.400 ;
        RECT  18.240 2.025 18.500 3.055 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.810 6.010 2.085 ;
        RECT  5.645 1.700 5.855 2.085 ;
        RECT  5.595 1.700 5.645 1.860 ;
        RECT  5.435 1.595 5.595 1.860 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.675 1.290 4.095 1.625 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 1.290 8.155 1.580 ;
        RECT  7.880 1.420 7.945 1.580 ;
        RECT  7.720 1.420 7.880 1.815 ;
        END
        ANTENNAGATEAREA     0.2366 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.195 -0.250 19.320 0.250 ;
        RECT  18.935 -0.250 19.195 1.095 ;
        RECT  18.145 -0.250 18.935 0.250 ;
        RECT  17.885 -0.250 18.145 0.565 ;
        RECT  17.065 -0.250 17.885 0.250 ;
        RECT  16.805 -0.250 17.065 0.405 ;
        RECT  16.260 -0.250 16.805 0.250 ;
        RECT  16.000 -0.250 16.260 0.405 ;
        RECT  13.270 -0.250 16.000 0.250 ;
        RECT  13.010 -0.250 13.270 0.960 ;
        RECT  12.200 -0.250 13.010 0.250 ;
        RECT  12.040 -0.250 12.200 1.295 ;
        RECT  10.430 -0.250 12.040 0.250 ;
        RECT  10.170 -0.250 10.430 0.950 ;
        RECT  9.100 -0.250 10.170 0.250 ;
        RECT  9.100 1.170 9.240 1.330 ;
        RECT  8.940 -0.250 9.100 1.330 ;
        RECT  8.300 -0.250 8.940 0.250 ;
        RECT  8.040 -0.250 8.300 0.405 ;
        RECT  5.870 -0.250 8.040 0.250 ;
        RECT  5.610 -0.250 5.870 0.405 ;
        RECT  3.925 -0.250 5.610 0.250 ;
        RECT  3.665 -0.250 3.925 0.405 ;
        RECT  1.525 -0.250 3.665 0.250 ;
        RECT  1.265 -0.250 1.525 0.405 ;
        RECT  0.385 -0.250 1.265 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.010 3.440 19.320 3.940 ;
        RECT  18.750 2.595 19.010 3.940 ;
        RECT  17.990 3.440 18.750 3.940 ;
        RECT  17.730 2.935 17.990 3.940 ;
        RECT  16.925 3.440 17.730 3.940 ;
        RECT  16.665 3.285 16.925 3.940 ;
        RECT  16.080 3.440 16.665 3.940 ;
        RECT  15.820 3.285 16.080 3.940 ;
        RECT  12.100 3.440 15.820 3.940 ;
        RECT  11.840 3.285 12.100 3.940 ;
        RECT  10.945 3.440 11.840 3.940 ;
        RECT  10.685 3.285 10.945 3.940 ;
        RECT  8.175 3.440 10.685 3.940 ;
        RECT  7.915 3.115 8.175 3.940 ;
        RECT  5.820 3.440 7.915 3.940 ;
        RECT  5.560 3.065 5.820 3.940 ;
        RECT  4.045 3.440 5.560 3.940 ;
        RECT  3.785 3.065 4.045 3.940 ;
        RECT  1.245 3.440 3.785 3.940 ;
        RECT  0.985 3.285 1.245 3.940 ;
        RECT  0.000 3.440 0.985 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.945 1.585 18.330 1.845 ;
        RECT  17.785 0.745 17.945 2.750 ;
        RECT  16.610 0.745 17.785 0.905 ;
        RECT  16.520 2.590 17.785 2.750 ;
        RECT  16.270 1.495 16.830 1.755 ;
        RECT  16.450 0.745 16.610 1.105 ;
        RECT  16.260 2.315 16.520 2.915 ;
        RECT  16.110 0.605 16.270 1.755 ;
        RECT  15.930 2.315 16.260 2.475 ;
        RECT  15.310 0.605 16.110 0.765 ;
        RECT  15.770 1.525 15.930 3.105 ;
        RECT  15.640 2.945 15.770 3.105 ;
        RECT  15.480 2.945 15.640 3.185 ;
        RECT  15.430 0.955 15.590 2.765 ;
        RECT  13.330 3.025 15.480 3.185 ;
        RECT  15.360 0.955 15.430 1.215 ;
        RECT  15.300 2.605 15.430 2.765 ;
        RECT  15.180 0.605 15.310 0.775 ;
        RECT  15.140 2.605 15.300 2.845 ;
        RECT  15.020 0.605 15.180 2.425 ;
        RECT  13.670 2.685 15.140 2.845 ;
        RECT  14.290 0.605 15.020 0.765 ;
        RECT  14.980 2.165 15.020 2.425 ;
        RECT  14.960 2.265 14.980 2.425 ;
        RECT  14.800 2.265 14.960 2.505 ;
        RECT  14.110 2.345 14.800 2.505 ;
        RECT  14.590 0.945 14.750 1.295 ;
        RECT  14.360 1.925 14.620 2.165 ;
        RECT  13.780 1.135 14.590 1.295 ;
        RECT  13.715 1.925 14.360 2.085 ;
        RECT  14.030 0.605 14.290 0.915 ;
        RECT  13.850 2.265 14.110 2.505 ;
        RECT  13.715 0.695 13.780 1.295 ;
        RECT  13.600 0.695 13.715 2.085 ;
        RECT  13.510 2.605 13.670 2.845 ;
        RECT  13.555 0.695 13.600 2.420 ;
        RECT  13.520 0.695 13.555 1.300 ;
        RECT  13.340 1.925 13.555 2.420 ;
        RECT  12.760 1.140 13.520 1.300 ;
        RECT  10.165 2.605 13.510 2.765 ;
        RECT  12.095 1.480 13.375 1.740 ;
        RECT  12.650 1.925 13.340 2.085 ;
        RECT  13.170 2.945 13.330 3.185 ;
        RECT  10.505 2.945 13.170 3.105 ;
        RECT  12.500 0.695 12.760 1.300 ;
        RECT  12.490 1.925 12.650 2.420 ;
        RECT  12.390 2.160 12.490 2.420 ;
        RECT  11.860 1.480 12.095 1.640 ;
        RECT  11.700 0.695 11.860 1.640 ;
        RECT  11.170 0.695 11.700 0.855 ;
        RECT  11.530 1.820 11.690 2.420 ;
        RECT  11.520 1.820 11.530 1.980 ;
        RECT  11.430 2.160 11.530 2.420 ;
        RECT  11.360 1.035 11.520 1.980 ;
        RECT  11.350 1.405 11.360 1.665 ;
        RECT  11.170 2.160 11.180 2.320 ;
        RECT  11.010 0.690 11.170 2.320 ;
        RECT  10.690 0.690 11.010 0.950 ;
        RECT  10.265 2.160 11.010 2.320 ;
        RECT  10.665 1.130 10.825 1.930 ;
        RECT  9.830 1.130 10.665 1.390 ;
        RECT  10.345 2.945 10.505 3.150 ;
        RECT  9.145 2.990 10.345 3.150 ;
        RECT  10.105 1.610 10.265 2.320 ;
        RECT  10.005 2.605 10.165 2.810 ;
        RECT  10.005 1.610 10.105 1.870 ;
        RECT  9.485 2.650 10.005 2.810 ;
        RECT  9.825 0.555 9.830 1.390 ;
        RECT  9.670 0.555 9.825 2.440 ;
        RECT  9.550 0.555 9.670 0.715 ;
        RECT  9.665 1.230 9.670 2.440 ;
        RECT  9.290 0.455 9.550 0.715 ;
        RECT  9.325 1.540 9.485 2.810 ;
        RECT  8.510 1.540 9.325 1.700 ;
        RECT  8.985 2.435 9.145 3.150 ;
        RECT  7.240 2.435 8.985 2.595 ;
        RECT  8.645 2.775 8.805 3.220 ;
        RECT  7.695 2.775 8.645 2.935 ;
        RECT  8.495 0.950 8.510 1.700 ;
        RECT  8.335 0.950 8.495 2.255 ;
        RECT  7.795 0.950 8.335 1.110 ;
        RECT  7.580 2.095 8.335 2.255 ;
        RECT  7.760 0.950 7.795 1.190 ;
        RECT  7.500 0.640 7.760 1.190 ;
        RECT  7.535 2.775 7.695 3.220 ;
        RECT  7.420 1.995 7.580 2.255 ;
        RECT  6.165 3.060 7.535 3.220 ;
        RECT  7.080 0.435 7.240 2.880 ;
        RECT  6.980 0.435 7.080 0.595 ;
        RECT  6.840 2.720 7.080 2.880 ;
        RECT  6.740 0.935 6.900 2.540 ;
        RECT  6.610 0.935 6.740 1.200 ;
        RECT  6.505 2.380 6.740 2.540 ;
        RECT  6.425 1.375 6.560 2.200 ;
        RECT  6.345 2.380 6.505 2.795 ;
        RECT  6.400 0.430 6.425 2.200 ;
        RECT  6.265 0.430 6.400 1.535 ;
        RECT  6.215 2.040 6.400 2.200 ;
        RECT  4.905 2.380 6.345 2.540 ;
        RECT  6.120 0.430 6.265 0.765 ;
        RECT  6.005 2.725 6.165 3.220 ;
        RECT  5.305 0.605 6.120 0.765 ;
        RECT  5.920 1.255 6.080 1.520 ;
        RECT  3.510 2.725 6.005 2.885 ;
        RECT  5.440 1.255 5.920 1.415 ;
        RECT  5.245 2.040 5.465 2.200 ;
        RECT  5.245 1.035 5.440 1.415 ;
        RECT  5.045 0.520 5.305 0.780 ;
        RECT  5.085 1.035 5.245 2.200 ;
        RECT  4.955 1.620 5.085 1.880 ;
        RECT  4.775 2.065 4.905 2.540 ;
        RECT  4.775 1.035 4.875 1.295 ;
        RECT  4.745 0.600 4.775 2.540 ;
        RECT  4.615 0.600 4.745 2.365 ;
        RECT  3.235 0.600 4.615 0.760 ;
        RECT  4.275 0.950 4.435 2.320 ;
        RECT  4.095 0.950 4.275 1.110 ;
        RECT  4.235 2.055 4.275 2.320 ;
        RECT  3.350 2.725 3.510 3.015 ;
        RECT  3.295 2.005 3.465 2.165 ;
        RECT  2.615 2.855 3.350 3.015 ;
        RECT  3.135 1.035 3.295 2.165 ;
        RECT  2.955 0.575 3.235 0.760 ;
        RECT  2.955 2.515 3.155 2.675 ;
        RECT  2.795 0.575 2.955 2.675 ;
        RECT  2.455 0.525 2.615 3.015 ;
        RECT  2.295 2.075 2.455 2.335 ;
        RECT  2.115 0.540 2.275 1.835 ;
        RECT  1.595 2.535 2.180 2.695 ;
        RECT  1.825 0.540 2.115 0.700 ;
        RECT  1.935 1.675 2.115 1.835 ;
        RECT  1.790 2.945 2.050 3.245 ;
        RECT  1.775 1.675 1.935 2.330 ;
        RECT  0.385 2.945 1.790 3.105 ;
        RECT  1.435 1.360 1.595 2.695 ;
        RECT  1.015 1.360 1.435 1.520 ;
        RECT  0.725 2.535 1.435 2.695 ;
        RECT  0.855 1.035 1.015 1.520 ;
        RECT  0.695 0.505 0.955 0.765 ;
        RECT  0.565 2.075 0.725 2.695 ;
        RECT  0.675 0.605 0.695 0.765 ;
        RECT  0.515 0.605 0.675 1.510 ;
        RECT  0.455 2.075 0.565 2.335 ;
        RECT  0.275 1.350 0.515 1.510 ;
        RECT  0.275 2.655 0.385 3.105 ;
        RECT  0.115 1.350 0.275 3.105 ;
    END
END SEDFFTRX4

MACRO SEDFFTRX2
    CLASS CORE ;
    FOREIGN SEDFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.775 1.010 1.935 1.495 ;
        RECT  1.715 1.010 1.775 1.170 ;
        RECT  1.505 0.880 1.715 1.170 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.910 1.700 1.255 2.080 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 0.635 0.335 1.170 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.915 2.145 16.965 2.405 ;
        RECT  16.685 0.820 16.915 2.405 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.235 0.690 18.275 1.500 ;
        RECT  18.090 0.600 18.235 1.500 ;
        RECT  17.985 0.600 18.090 1.580 ;
        RECT  17.975 0.600 17.985 3.100 ;
        RECT  17.825 1.340 17.975 3.100 ;
        RECT  17.725 2.110 17.825 3.100 ;
        RECT  17.605 2.110 17.725 2.585 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.810 6.010 2.085 ;
        RECT  5.645 1.670 5.855 2.085 ;
        RECT  5.425 1.670 5.645 1.830 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.675 1.290 4.095 1.625 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 1.290 8.155 1.580 ;
        RECT  7.925 1.420 7.945 1.580 ;
        RECT  7.765 1.420 7.925 1.815 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.695 -0.250 18.400 0.250 ;
        RECT  17.435 -0.250 17.695 1.135 ;
        RECT  15.905 -0.250 17.435 0.250 ;
        RECT  15.645 -0.250 15.905 0.405 ;
        RECT  13.285 -0.250 15.645 0.250 ;
        RECT  13.025 -0.250 13.285 0.785 ;
        RECT  12.180 -0.250 13.025 0.250 ;
        RECT  12.020 -0.250 12.180 1.130 ;
        RECT  10.420 -0.250 12.020 0.250 ;
        RECT  10.160 -0.250 10.420 0.950 ;
        RECT  9.100 -0.250 10.160 0.250 ;
        RECT  9.100 1.170 9.225 1.330 ;
        RECT  8.940 -0.250 9.100 1.330 ;
        RECT  8.275 -0.250 8.940 0.250 ;
        RECT  8.015 -0.250 8.275 0.405 ;
        RECT  5.870 -0.250 8.015 0.250 ;
        RECT  5.610 -0.250 5.870 0.405 ;
        RECT  3.925 -0.250 5.610 0.250 ;
        RECT  3.665 -0.250 3.925 0.405 ;
        RECT  1.525 -0.250 3.665 0.250 ;
        RECT  1.265 -0.250 1.525 0.405 ;
        RECT  0.385 -0.250 1.265 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.475 3.440 18.400 3.940 ;
        RECT  17.215 2.935 17.475 3.940 ;
        RECT  15.905 3.440 17.215 3.940 ;
        RECT  15.645 3.285 15.905 3.940 ;
        RECT  13.030 3.440 15.645 3.940 ;
        RECT  12.770 3.285 13.030 3.940 ;
        RECT  12.080 3.440 12.770 3.940 ;
        RECT  11.820 3.285 12.080 3.940 ;
        RECT  10.945 3.440 11.820 3.940 ;
        RECT  10.685 3.285 10.945 3.940 ;
        RECT  8.175 3.440 10.685 3.940 ;
        RECT  7.915 3.115 8.175 3.940 ;
        RECT  5.825 3.440 7.915 3.940 ;
        RECT  5.565 3.065 5.825 3.940 ;
        RECT  4.045 3.440 5.565 3.940 ;
        RECT  3.785 3.065 4.045 3.940 ;
        RECT  1.245 3.440 3.785 3.940 ;
        RECT  0.985 3.285 1.245 3.940 ;
        RECT  0.000 3.440 0.985 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.305 1.585 17.645 1.845 ;
        RECT  17.255 1.585 17.305 2.755 ;
        RECT  17.145 0.475 17.255 2.755 ;
        RECT  17.095 0.475 17.145 1.745 ;
        RECT  16.455 2.595 17.145 2.755 ;
        RECT  16.455 0.475 17.095 0.635 ;
        RECT  16.295 0.475 16.455 1.095 ;
        RECT  16.195 2.190 16.455 3.105 ;
        RECT  16.195 0.835 16.295 1.095 ;
        RECT  16.100 1.635 16.285 1.895 ;
        RECT  15.755 2.945 16.195 3.105 ;
        RECT  15.940 1.280 16.100 1.895 ;
        RECT  15.650 1.280 15.940 1.440 ;
        RECT  15.595 1.620 15.755 3.105 ;
        RECT  15.490 0.770 15.650 1.440 ;
        RECT  10.505 2.945 15.595 3.105 ;
        RECT  15.120 0.770 15.490 0.930 ;
        RECT  15.275 1.680 15.390 2.765 ;
        RECT  15.230 1.330 15.275 2.765 ;
        RECT  15.115 1.330 15.230 1.840 ;
        RECT  11.860 2.605 15.230 2.765 ;
        RECT  14.930 0.770 15.120 1.150 ;
        RECT  14.930 2.020 15.050 2.280 ;
        RECT  14.770 0.770 14.930 2.425 ;
        RECT  14.210 0.845 14.770 1.005 ;
        RECT  13.790 2.265 14.770 2.425 ;
        RECT  14.595 0.430 14.760 0.590 ;
        RECT  14.435 0.430 14.595 0.665 ;
        RECT  13.540 1.925 14.590 2.085 ;
        RECT  13.650 0.505 14.435 0.665 ;
        RECT  13.950 0.845 14.210 1.105 ;
        RECT  13.490 0.505 13.650 1.295 ;
        RECT  13.280 1.925 13.540 2.215 ;
        RECT  13.390 1.035 13.490 1.295 ;
        RECT  12.790 1.035 13.390 1.200 ;
        RECT  12.790 1.925 13.280 2.090 ;
        RECT  12.630 1.035 12.790 2.090 ;
        RECT  12.480 1.035 12.630 1.295 ;
        RECT  12.370 1.930 12.630 2.215 ;
        RECT  12.165 1.480 12.425 1.740 ;
        RECT  11.840 1.480 12.165 1.640 ;
        RECT  11.650 2.600 11.860 2.765 ;
        RECT  11.680 0.690 11.840 1.640 ;
        RECT  11.430 1.915 11.690 2.215 ;
        RECT  10.930 0.690 11.680 0.850 ;
        RECT  10.165 2.600 11.650 2.760 ;
        RECT  11.400 1.035 11.500 1.295 ;
        RECT  11.400 1.915 11.430 2.075 ;
        RECT  11.240 1.035 11.400 2.075 ;
        RECT  11.050 1.410 11.240 1.670 ;
        RECT  10.870 2.260 11.180 2.420 ;
        RECT  10.870 0.690 10.930 0.950 ;
        RECT  10.710 0.690 10.870 2.420 ;
        RECT  10.670 0.690 10.710 0.950 ;
        RECT  10.275 2.260 10.710 2.420 ;
        RECT  9.830 1.130 10.530 1.390 ;
        RECT  10.345 2.945 10.505 3.150 ;
        RECT  10.275 1.610 10.395 1.870 ;
        RECT  9.145 2.990 10.345 3.150 ;
        RECT  10.115 1.610 10.275 2.420 ;
        RECT  10.005 2.600 10.165 2.810 ;
        RECT  9.485 2.650 10.005 2.810 ;
        RECT  9.825 0.555 9.830 1.390 ;
        RECT  9.670 0.555 9.825 2.440 ;
        RECT  9.540 0.555 9.670 0.715 ;
        RECT  9.665 1.230 9.670 2.440 ;
        RECT  9.280 0.455 9.540 0.715 ;
        RECT  9.325 1.540 9.485 2.810 ;
        RECT  8.510 1.540 9.325 1.700 ;
        RECT  8.985 2.435 9.145 3.150 ;
        RECT  7.355 2.435 8.985 2.595 ;
        RECT  8.645 2.775 8.805 3.220 ;
        RECT  7.695 2.775 8.645 2.935 ;
        RECT  8.495 0.950 8.510 1.700 ;
        RECT  8.335 0.950 8.495 2.255 ;
        RECT  7.795 0.950 8.335 1.110 ;
        RECT  7.695 2.095 8.335 2.255 ;
        RECT  7.610 0.475 7.795 1.110 ;
        RECT  7.535 1.995 7.695 2.255 ;
        RECT  7.535 2.775 7.695 3.220 ;
        RECT  7.505 0.475 7.610 0.635 ;
        RECT  6.165 3.060 7.535 3.220 ;
        RECT  7.195 0.935 7.355 2.880 ;
        RECT  6.840 2.720 7.195 2.880 ;
        RECT  6.855 0.530 7.015 2.540 ;
        RECT  6.810 0.530 6.855 0.690 ;
        RECT  6.505 2.380 6.855 2.540 ;
        RECT  6.550 0.430 6.810 0.690 ;
        RECT  6.535 1.620 6.675 1.885 ;
        RECT  6.375 0.990 6.535 2.200 ;
        RECT  6.345 2.380 6.505 2.795 ;
        RECT  6.035 0.990 6.375 1.150 ;
        RECT  6.215 2.040 6.375 2.200 ;
        RECT  4.905 2.380 6.345 2.540 ;
        RECT  6.035 1.330 6.195 1.590 ;
        RECT  6.005 2.720 6.165 3.220 ;
        RECT  5.875 0.605 6.035 1.150 ;
        RECT  5.440 1.330 6.035 1.490 ;
        RECT  3.510 2.720 6.005 2.880 ;
        RECT  5.295 0.605 5.875 0.765 ;
        RECT  5.245 2.040 5.465 2.200 ;
        RECT  5.245 1.035 5.440 1.490 ;
        RECT  5.035 0.595 5.295 0.855 ;
        RECT  5.180 1.035 5.245 2.200 ;
        RECT  5.085 1.330 5.180 2.200 ;
        RECT  4.955 1.620 5.085 1.880 ;
        RECT  4.775 2.065 4.905 2.540 ;
        RECT  4.775 1.035 4.875 1.295 ;
        RECT  4.745 0.600 4.775 2.540 ;
        RECT  4.615 0.600 4.745 2.365 ;
        RECT  3.235 0.600 4.615 0.760 ;
        RECT  4.275 0.950 4.435 2.320 ;
        RECT  4.095 0.950 4.275 1.110 ;
        RECT  4.235 2.055 4.275 2.320 ;
        RECT  3.350 2.720 3.510 3.015 ;
        RECT  3.295 2.005 3.465 2.165 ;
        RECT  2.615 2.855 3.350 3.015 ;
        RECT  3.135 1.035 3.295 2.165 ;
        RECT  2.955 0.575 3.235 0.760 ;
        RECT  2.955 2.515 3.155 2.675 ;
        RECT  2.795 0.575 2.955 2.675 ;
        RECT  2.455 0.525 2.615 3.015 ;
        RECT  2.295 2.065 2.455 2.325 ;
        RECT  2.115 0.540 2.275 1.835 ;
        RECT  1.920 2.505 2.180 2.765 ;
        RECT  1.825 0.540 2.115 0.700 ;
        RECT  1.935 1.675 2.115 1.835 ;
        RECT  1.790 2.945 2.050 3.245 ;
        RECT  1.775 1.675 1.935 2.325 ;
        RECT  1.595 2.605 1.920 2.765 ;
        RECT  0.385 2.945 1.790 3.105 ;
        RECT  1.435 1.360 1.595 2.765 ;
        RECT  1.015 1.360 1.435 1.520 ;
        RECT  0.725 2.605 1.435 2.765 ;
        RECT  0.855 1.035 1.015 1.520 ;
        RECT  0.675 0.555 0.955 0.715 ;
        RECT  0.565 2.075 0.725 2.765 ;
        RECT  0.515 0.555 0.675 1.510 ;
        RECT  0.455 2.075 0.565 2.335 ;
        RECT  0.275 1.350 0.515 1.510 ;
        RECT  0.275 2.655 0.385 3.105 ;
        RECT  0.115 1.350 0.275 3.105 ;
    END
END SEDFFTRX2

MACRO SEDFFTRX1
    CLASS CORE ;
    FOREIGN SEDFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.100 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.010 1.825 1.495 ;
        RECT  1.665 0.880 1.715 1.495 ;
        RECT  1.505 0.880 1.665 1.170 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.700 1.115 2.035 ;
        RECT  0.585 1.700 0.905 1.990 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 0.585 0.335 1.170 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.975 0.975 15.055 2.215 ;
        RECT  14.845 0.975 14.975 2.595 ;
        RECT  14.695 0.975 14.845 1.235 ;
        RECT  14.715 1.995 14.845 2.595 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.925 0.975 15.975 2.175 ;
        RECT  15.765 0.975 15.925 2.595 ;
        RECT  15.645 0.975 15.765 1.235 ;
        RECT  15.665 1.995 15.765 2.595 ;
        END
        ANTENNADIFFAREA     0.3538 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.775 6.035 2.200 ;
        RECT  5.675 1.700 5.855 2.200 ;
        RECT  5.640 1.670 5.675 2.200 ;
        RECT  5.415 1.670 5.640 1.860 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.370 4.095 1.990 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 1.290 8.155 1.580 ;
        RECT  7.755 1.420 7.945 1.580 ;
        RECT  7.495 1.405 7.755 1.665 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.355 -0.250 16.100 0.250 ;
        RECT  15.095 -0.250 15.355 0.405 ;
        RECT  14.085 -0.250 15.095 0.250 ;
        RECT  13.825 -0.250 14.085 0.405 ;
        RECT  12.065 -0.250 13.825 0.250 ;
        RECT  11.805 -0.250 12.065 0.610 ;
        RECT  10.475 -0.250 11.805 0.250 ;
        RECT  10.215 -0.250 10.475 0.950 ;
        RECT  9.065 -0.250 10.215 0.250 ;
        RECT  8.805 -0.250 9.065 1.385 ;
        RECT  8.125 -0.250 8.805 0.250 ;
        RECT  7.865 -0.250 8.125 0.745 ;
        RECT  5.875 -0.250 7.865 0.250 ;
        RECT  5.615 -0.250 5.875 0.405 ;
        RECT  3.785 -0.250 5.615 0.250 ;
        RECT  3.525 -0.250 3.785 0.405 ;
        RECT  1.525 -0.250 3.525 0.250 ;
        RECT  1.265 -0.250 1.525 0.405 ;
        RECT  0.385 -0.250 1.265 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.375 3.440 16.100 3.940 ;
        RECT  15.115 3.285 15.375 3.940 ;
        RECT  13.975 3.440 15.115 3.940 ;
        RECT  13.715 3.285 13.975 3.940 ;
        RECT  12.135 3.440 13.715 3.940 ;
        RECT  11.875 3.285 12.135 3.940 ;
        RECT  10.765 3.440 11.875 3.940 ;
        RECT  10.505 3.285 10.765 3.940 ;
        RECT  8.175 3.440 10.505 3.940 ;
        RECT  7.915 3.115 8.175 3.940 ;
        RECT  5.775 3.440 7.915 3.940 ;
        RECT  5.515 3.115 5.775 3.940 ;
        RECT  4.035 3.440 5.515 3.940 ;
        RECT  3.775 3.115 4.035 3.940 ;
        RECT  1.215 3.440 3.775 3.940 ;
        RECT  0.955 3.285 1.215 3.940 ;
        RECT  0.000 3.440 0.955 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.465 1.475 15.585 1.735 ;
        RECT  15.305 0.585 15.465 3.005 ;
        RECT  14.595 0.585 15.305 0.745 ;
        RECT  14.615 2.845 15.305 3.005 ;
        RECT  14.355 2.845 14.615 3.105 ;
        RECT  14.335 0.430 14.595 0.745 ;
        RECT  14.395 1.495 14.495 1.755 ;
        RECT  14.235 0.985 14.395 1.755 ;
        RECT  13.875 2.945 14.355 3.105 ;
        RECT  13.685 0.985 14.235 1.145 ;
        RECT  13.715 1.325 13.875 3.105 ;
        RECT  13.615 1.325 13.715 1.585 ;
        RECT  10.315 2.945 13.715 3.105 ;
        RECT  13.525 0.615 13.685 1.145 ;
        RECT  13.005 0.615 13.525 0.775 ;
        RECT  13.355 1.765 13.515 2.765 ;
        RECT  13.345 1.765 13.355 1.925 ;
        RECT  13.225 2.600 13.355 2.765 ;
        RECT  13.185 0.955 13.345 1.925 ;
        RECT  11.905 2.600 13.225 2.760 ;
        RECT  13.005 2.150 13.175 2.410 ;
        RECT  12.845 0.615 13.005 2.410 ;
        RECT  12.505 0.685 12.665 2.420 ;
        RECT  12.355 0.685 12.505 1.235 ;
        RECT  12.055 1.445 12.315 1.705 ;
        RECT  11.975 1.445 12.055 1.605 ;
        RECT  11.815 0.790 11.975 1.605 ;
        RECT  11.645 2.590 11.905 2.760 ;
        RECT  11.045 0.790 11.815 0.950 ;
        RECT  11.585 2.200 11.705 2.360 ;
        RECT  9.970 2.600 11.645 2.760 ;
        RECT  11.585 1.130 11.635 1.290 ;
        RECT  11.425 1.130 11.585 2.360 ;
        RECT  11.375 1.130 11.425 1.290 ;
        RECT  11.155 1.470 11.425 1.730 ;
        RECT  10.975 2.260 11.195 2.420 ;
        RECT  10.975 0.690 11.045 0.950 ;
        RECT  10.815 0.690 10.975 2.420 ;
        RECT  10.785 0.690 10.815 0.950 ;
        RECT  10.275 1.710 10.815 1.870 ;
        RECT  9.835 1.130 10.635 1.390 ;
        RECT  10.155 2.945 10.315 3.150 ;
        RECT  10.015 1.610 10.275 1.870 ;
        RECT  9.155 2.990 10.155 3.150 ;
        RECT  9.710 2.600 9.970 2.810 ;
        RECT  9.675 0.705 9.835 2.345 ;
        RECT  9.495 2.600 9.710 2.760 ;
        RECT  9.595 0.705 9.675 0.865 ;
        RECT  9.335 0.540 9.595 0.865 ;
        RECT  9.335 1.045 9.495 2.760 ;
        RECT  9.245 1.045 9.335 1.305 ;
        RECT  8.495 1.795 9.335 1.955 ;
        RECT  8.995 2.140 9.155 3.150 ;
        RECT  8.435 2.140 8.995 2.300 ;
        RECT  8.655 2.545 8.815 2.935 ;
        RECT  7.695 2.775 8.655 2.935 ;
        RECT  8.335 0.950 8.495 1.955 ;
        RECT  8.275 2.140 8.435 2.590 ;
        RECT  7.685 0.950 8.335 1.110 ;
        RECT  8.095 1.795 8.335 1.955 ;
        RECT  7.355 2.430 8.275 2.590 ;
        RECT  7.935 1.795 8.095 2.060 ;
        RECT  7.695 1.900 7.935 2.060 ;
        RECT  7.535 1.900 7.695 2.250 ;
        RECT  7.535 2.775 7.695 3.220 ;
        RECT  7.525 0.585 7.685 1.110 ;
        RECT  6.115 3.060 7.535 3.220 ;
        RECT  7.405 0.585 7.525 0.745 ;
        RECT  7.145 0.495 7.405 0.745 ;
        RECT  7.315 2.430 7.355 2.880 ;
        RECT  7.155 1.035 7.315 2.880 ;
        RECT  6.805 2.720 7.155 2.880 ;
        RECT  6.895 1.030 6.975 2.540 ;
        RECT  6.815 0.430 6.895 2.540 ;
        RECT  6.735 0.430 6.815 1.190 ;
        RECT  6.555 2.380 6.815 2.540 ;
        RECT  6.635 0.430 6.735 0.590 ;
        RECT  6.535 1.620 6.635 1.880 ;
        RECT  6.395 2.380 6.555 2.880 ;
        RECT  6.395 0.770 6.535 2.200 ;
        RECT  6.375 0.470 6.395 2.200 ;
        RECT  6.295 2.435 6.395 2.880 ;
        RECT  6.235 0.470 6.375 0.930 ;
        RECT  6.215 2.040 6.375 2.200 ;
        RECT  4.895 2.435 6.295 2.595 ;
        RECT  6.125 0.470 6.235 0.765 ;
        RECT  5.895 1.260 6.155 1.520 ;
        RECT  5.245 0.605 6.125 0.765 ;
        RECT  5.955 2.775 6.115 3.220 ;
        RECT  3.395 2.775 5.955 2.935 ;
        RECT  5.445 1.330 5.895 1.490 ;
        RECT  5.235 2.040 5.455 2.200 ;
        RECT  5.235 0.955 5.445 1.490 ;
        RECT  4.985 0.515 5.245 0.775 ;
        RECT  5.185 0.955 5.235 2.200 ;
        RECT  5.075 1.330 5.185 2.200 ;
        RECT  4.985 1.620 5.075 1.880 ;
        RECT  4.805 0.965 4.935 1.125 ;
        RECT  4.805 2.265 4.895 2.595 ;
        RECT  4.645 0.585 4.805 2.595 ;
        RECT  3.215 0.585 4.645 0.745 ;
        RECT  4.275 0.925 4.435 2.545 ;
        RECT  4.105 0.925 4.275 1.185 ;
        RECT  4.175 2.285 4.275 2.545 ;
        RECT  3.295 2.195 3.465 2.455 ;
        RECT  3.235 2.775 3.395 3.065 ;
        RECT  3.135 1.035 3.295 2.455 ;
        RECT  2.515 2.905 3.235 3.065 ;
        RECT  2.955 0.575 3.215 0.745 ;
        RECT  2.795 0.575 2.955 2.725 ;
        RECT  2.695 2.465 2.795 2.725 ;
        RECT  2.515 0.640 2.595 2.250 ;
        RECT  2.435 0.640 2.515 3.065 ;
        RECT  2.355 2.090 2.435 3.065 ;
        RECT  2.155 2.090 2.355 2.350 ;
        RECT  2.005 0.540 2.165 1.835 ;
        RECT  1.815 0.540 2.005 0.700 ;
        RECT  1.795 1.675 2.005 1.835 ;
        RECT  1.715 2.505 1.975 2.765 ;
        RECT  1.705 2.945 1.965 3.245 ;
        RECT  1.635 1.675 1.795 2.305 ;
        RECT  1.455 2.605 1.715 2.765 ;
        RECT  0.385 2.945 1.705 3.105 ;
        RECT  1.295 1.360 1.455 2.765 ;
        RECT  1.015 1.360 1.295 1.520 ;
        RECT  0.725 2.605 1.295 2.765 ;
        RECT  0.855 1.035 1.015 1.520 ;
        RECT  0.695 0.555 0.955 0.855 ;
        RECT  0.565 2.170 0.725 2.765 ;
        RECT  0.675 0.695 0.695 0.855 ;
        RECT  0.515 0.695 0.675 1.510 ;
        RECT  0.465 2.170 0.565 2.335 ;
        RECT  0.285 1.350 0.515 1.510 ;
        RECT  0.285 2.700 0.385 3.105 ;
        RECT  0.125 1.350 0.285 3.105 ;
    END
END SEDFFTRX1

MACRO SEDFFTRXL
    CLASS CORE ;
    FOREIGN SEDFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.640 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.775 1.010 1.935 1.495 ;
        RECT  1.715 1.010 1.775 1.170 ;
        RECT  1.505 0.880 1.715 1.170 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.855 1.700 1.255 2.135 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.105 0.705 0.335 1.545 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.595 1.290 14.735 2.570 ;
        RECT  14.575 0.940 14.595 2.570 ;
        RECT  14.385 0.940 14.575 1.580 ;
        RECT  14.255 2.310 14.575 2.570 ;
        RECT  14.285 0.940 14.385 1.100 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.355 0.880 15.515 2.425 ;
        RECT  15.330 0.880 15.355 1.360 ;
        RECT  15.255 2.165 15.355 2.425 ;
        RECT  15.305 0.880 15.330 1.295 ;
        RECT  15.255 1.035 15.305 1.295 ;
        END
        ANTENNADIFFAREA     0.2312 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.775 6.035 2.200 ;
        RECT  5.640 1.670 5.855 2.200 ;
        RECT  5.415 1.670 5.640 1.860 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.380 4.085 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 1.290 8.155 1.580 ;
        RECT  7.825 1.420 7.945 1.580 ;
        RECT  7.665 1.420 7.825 1.685 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.055 -0.250 15.640 0.250 ;
        RECT  14.795 -0.250 15.055 0.405 ;
        RECT  13.965 -0.250 14.795 0.250 ;
        RECT  13.705 -0.250 13.965 0.405 ;
        RECT  12.265 -0.250 13.705 0.250 ;
        RECT  12.105 -0.250 12.265 0.785 ;
        RECT  10.475 -0.250 12.105 0.250 ;
        RECT  10.215 -0.250 10.475 0.950 ;
        RECT  8.835 -0.250 10.215 0.250 ;
        RECT  8.835 1.125 8.995 1.385 ;
        RECT  8.675 -0.250 8.835 1.385 ;
        RECT  8.125 -0.250 8.675 0.250 ;
        RECT  7.865 -0.250 8.125 0.405 ;
        RECT  6.065 -0.250 7.865 0.250 ;
        RECT  5.805 -0.250 6.065 0.405 ;
        RECT  3.860 -0.250 5.805 0.250 ;
        RECT  3.600 -0.250 3.860 0.405 ;
        RECT  1.525 -0.250 3.600 0.250 ;
        RECT  1.265 -0.250 1.525 0.405 ;
        RECT  0.385 -0.250 1.265 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.055 3.440 15.640 3.940 ;
        RECT  14.795 3.285 15.055 3.940 ;
        RECT  13.975 3.440 14.795 3.940 ;
        RECT  13.715 3.285 13.975 3.940 ;
        RECT  12.170 3.440 13.715 3.940 ;
        RECT  11.910 3.285 12.170 3.940 ;
        RECT  10.765 3.440 11.910 3.940 ;
        RECT  10.505 3.285 10.765 3.940 ;
        RECT  8.175 3.440 10.505 3.940 ;
        RECT  7.915 3.115 8.175 3.940 ;
        RECT  5.770 3.440 7.915 3.940 ;
        RECT  5.510 3.115 5.770 3.940 ;
        RECT  4.005 3.440 5.510 3.940 ;
        RECT  3.745 3.115 4.005 3.940 ;
        RECT  1.095 3.440 3.745 3.940 ;
        RECT  0.835 3.285 1.095 3.940 ;
        RECT  0.000 3.440 0.835 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.075 1.635 15.175 1.895 ;
        RECT  14.915 0.585 15.075 2.910 ;
        RECT  14.545 0.585 14.915 0.745 ;
        RECT  14.545 2.750 14.915 2.910 ;
        RECT  14.285 0.430 14.545 0.745 ;
        RECT  14.285 2.750 14.545 3.120 ;
        RECT  14.205 1.760 14.385 2.020 ;
        RECT  13.855 2.945 14.285 3.105 ;
        RECT  14.045 1.280 14.205 2.020 ;
        RECT  13.720 1.280 14.045 1.440 ;
        RECT  13.695 1.620 13.855 3.105 ;
        RECT  13.560 0.630 13.720 1.440 ;
        RECT  10.315 2.945 13.695 3.105 ;
        RECT  13.005 0.630 13.560 0.790 ;
        RECT  13.375 1.680 13.515 2.760 ;
        RECT  13.355 1.020 13.375 2.760 ;
        RECT  13.215 1.020 13.355 1.840 ;
        RECT  9.970 2.600 13.355 2.760 ;
        RECT  13.005 2.020 13.175 2.280 ;
        RECT  12.845 0.630 13.005 2.280 ;
        RECT  12.505 1.035 12.665 2.280 ;
        RECT  12.385 1.035 12.505 1.295 ;
        RECT  12.065 1.480 12.325 1.740 ;
        RECT  11.925 1.480 12.065 1.640 ;
        RECT  11.765 0.685 11.925 1.640 ;
        RECT  11.045 0.685 11.765 0.845 ;
        RECT  11.585 2.220 11.705 2.380 ;
        RECT  11.425 1.025 11.585 1.290 ;
        RECT  11.425 1.915 11.585 2.380 ;
        RECT  11.415 1.130 11.425 1.290 ;
        RECT  11.315 1.915 11.425 2.075 ;
        RECT  11.315 1.130 11.415 1.665 ;
        RECT  11.255 1.130 11.315 2.075 ;
        RECT  11.155 1.405 11.255 2.075 ;
        RECT  10.975 2.260 11.195 2.420 ;
        RECT  10.975 0.685 11.045 0.950 ;
        RECT  10.815 0.685 10.975 2.420 ;
        RECT  10.785 0.690 10.815 0.950 ;
        RECT  10.275 2.260 10.815 2.420 ;
        RECT  9.835 1.130 10.635 1.390 ;
        RECT  10.155 2.945 10.315 3.150 ;
        RECT  10.115 1.610 10.275 2.420 ;
        RECT  9.155 2.990 10.155 3.150 ;
        RECT  10.015 1.610 10.115 1.870 ;
        RECT  9.710 2.600 9.970 2.810 ;
        RECT  9.815 1.130 9.835 2.345 ;
        RECT  9.675 0.705 9.815 2.345 ;
        RECT  9.495 2.600 9.710 2.760 ;
        RECT  9.655 0.705 9.675 1.290 ;
        RECT  9.595 0.705 9.655 0.865 ;
        RECT  9.335 0.605 9.595 0.865 ;
        RECT  9.475 1.495 9.495 2.760 ;
        RECT  9.335 1.045 9.475 2.760 ;
        RECT  9.315 1.045 9.335 2.025 ;
        RECT  9.175 1.045 9.315 1.305 ;
        RECT  8.495 1.865 9.315 2.025 ;
        RECT  8.995 2.205 9.155 3.150 ;
        RECT  8.070 2.205 8.995 2.365 ;
        RECT  8.655 2.545 8.815 2.935 ;
        RECT  7.695 2.775 8.655 2.935 ;
        RECT  8.335 0.950 8.495 2.025 ;
        RECT  7.695 0.950 8.335 1.110 ;
        RECT  7.695 1.865 8.335 2.025 ;
        RECT  7.910 2.205 8.070 2.595 ;
        RECT  7.355 2.435 7.910 2.595 ;
        RECT  7.545 0.585 7.695 1.110 ;
        RECT  7.535 1.865 7.695 2.255 ;
        RECT  7.535 2.775 7.695 3.220 ;
        RECT  7.535 0.475 7.545 1.110 ;
        RECT  7.280 0.475 7.535 0.750 ;
        RECT  6.115 3.060 7.535 3.220 ;
        RECT  7.195 0.935 7.355 2.880 ;
        RECT  6.805 2.720 7.195 2.880 ;
        RECT  6.875 0.940 7.015 2.540 ;
        RECT  6.855 0.430 6.875 2.540 ;
        RECT  6.715 0.430 6.855 1.100 ;
        RECT  6.555 2.380 6.855 2.540 ;
        RECT  6.580 0.430 6.715 0.690 ;
        RECT  6.535 1.620 6.675 1.885 ;
        RECT  6.295 2.380 6.555 2.880 ;
        RECT  6.395 0.990 6.535 2.200 ;
        RECT  6.375 0.585 6.395 2.200 ;
        RECT  6.235 0.585 6.375 1.150 ;
        RECT  6.215 2.040 6.375 2.200 ;
        RECT  4.895 2.380 6.295 2.540 ;
        RECT  5.210 0.585 6.235 0.745 ;
        RECT  6.035 1.330 6.195 1.590 ;
        RECT  5.955 2.725 6.115 3.220 ;
        RECT  5.485 1.330 6.035 1.490 ;
        RECT  3.395 2.725 5.955 2.885 ;
        RECT  5.235 1.005 5.485 1.490 ;
        RECT  5.235 2.040 5.455 2.200 ;
        RECT  5.225 1.005 5.235 2.200 ;
        RECT  5.075 1.330 5.225 2.200 ;
        RECT  4.950 0.550 5.210 0.810 ;
        RECT  4.950 1.620 5.075 1.880 ;
        RECT  4.770 0.990 4.975 1.150 ;
        RECT  4.770 2.265 4.895 2.540 ;
        RECT  4.610 0.600 4.770 2.540 ;
        RECT  3.205 0.600 4.610 0.760 ;
        RECT  4.270 0.940 4.430 2.435 ;
        RECT  4.170 0.940 4.270 1.200 ;
        RECT  4.175 2.175 4.270 2.435 ;
        RECT  3.295 1.955 3.415 2.215 ;
        RECT  3.235 2.725 3.395 3.065 ;
        RECT  3.135 1.035 3.295 2.215 ;
        RECT  2.615 2.905 3.235 3.065 ;
        RECT  2.955 0.490 3.205 0.760 ;
        RECT  2.955 2.465 3.055 2.725 ;
        RECT  2.945 0.490 2.955 2.725 ;
        RECT  2.795 0.600 2.945 2.725 ;
        RECT  2.455 0.490 2.615 3.065 ;
        RECT  2.235 2.115 2.455 2.375 ;
        RECT  2.115 0.540 2.275 1.835 ;
        RECT  1.815 0.540 2.115 0.700 ;
        RECT  1.935 1.675 2.115 1.835 ;
        RECT  1.595 2.555 2.105 2.765 ;
        RECT  1.790 2.985 2.050 3.245 ;
        RECT  1.775 1.675 1.935 2.215 ;
        RECT  1.435 2.985 1.790 3.145 ;
        RECT  1.435 1.360 1.595 2.765 ;
        RECT  1.015 1.360 1.435 1.520 ;
        RECT  0.725 2.605 1.435 2.765 ;
        RECT  1.275 2.945 1.435 3.145 ;
        RECT  0.385 2.945 1.275 3.105 ;
        RECT  0.855 1.035 1.015 1.520 ;
        RECT  0.695 0.505 0.955 0.855 ;
        RECT  0.615 2.315 0.725 2.765 ;
        RECT  0.675 0.695 0.695 0.855 ;
        RECT  0.515 0.695 0.675 1.890 ;
        RECT  0.565 2.075 0.615 2.765 ;
        RECT  0.455 2.075 0.565 2.475 ;
        RECT  0.275 1.730 0.515 1.890 ;
        RECT  0.275 2.655 0.385 3.105 ;
        RECT  0.115 1.730 0.275 3.105 ;
    END
END SEDFFTRXL

MACRO SEDFFX4
    CLASS CORE ;
    FOREIGN SEDFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.100 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 1.655 2.640 1.990 ;
        END
        ANTENNAGATEAREA     0.1131 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.700 1.530 1.990 ;
        END
        ANTENNAGATEAREA     0.1807 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.505 1.515 15.515 2.585 ;
        RECT  15.455 0.920 15.505 2.585 ;
        RECT  15.440 0.920 15.455 3.030 ;
        RECT  15.305 0.590 15.440 3.030 ;
        RECT  15.180 0.590 15.305 1.190 ;
        RECT  15.195 2.090 15.305 3.030 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.425 1.700 14.435 2.400 ;
        RECT  14.420 0.810 14.425 2.400 ;
        RECT  14.265 0.590 14.420 2.400 ;
        RECT  14.160 0.590 14.265 1.190 ;
        RECT  13.925 1.700 14.265 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.650 0.525 3.050 ;
        RECT  0.265 2.520 0.335 3.050 ;
        RECT  0.125 2.520 0.265 2.810 ;
        END
        ANTENNAGATEAREA     0.1781 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.275 1.610 3.495 1.865 ;
        RECT  3.085 1.610 3.275 1.990 ;
        RECT  2.885 1.700 3.085 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 1.675 7.130 1.990 ;
        END
        ANTENNAGATEAREA     0.2340 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.950 -0.250 16.100 0.250 ;
        RECT  15.690 -0.250 15.950 1.190 ;
        RECT  14.930 -0.250 15.690 0.250 ;
        RECT  14.670 -0.250 14.930 1.190 ;
        RECT  13.910 -0.250 14.670 0.250 ;
        RECT  13.650 -0.250 13.910 1.190 ;
        RECT  12.760 -0.250 13.650 0.250 ;
        RECT  12.500 -0.250 12.760 1.210 ;
        RECT  10.745 -0.250 12.500 0.250 ;
        RECT  10.485 -0.250 10.745 0.885 ;
        RECT  9.070 -0.250 10.485 0.250 ;
        RECT  8.810 -0.250 9.070 0.955 ;
        RECT  7.390 -0.250 8.810 0.250 ;
        RECT  7.130 -0.250 7.390 0.405 ;
        RECT  6.430 -0.250 7.130 0.250 ;
        RECT  6.170 -0.250 6.430 0.405 ;
        RECT  2.550 -0.250 6.170 0.250 ;
        RECT  2.290 -0.250 2.550 0.665 ;
        RECT  0.965 -0.250 2.290 0.250 ;
        RECT  0.705 -0.250 0.965 0.795 ;
        RECT  0.000 -0.250 0.705 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.965 3.440 16.100 3.940 ;
        RECT  15.705 2.210 15.965 3.940 ;
        RECT  14.945 3.440 15.705 3.940 ;
        RECT  14.685 2.930 14.945 3.940 ;
        RECT  13.925 3.440 14.685 3.940 ;
        RECT  13.665 2.935 13.925 3.940 ;
        RECT  12.875 3.440 13.665 3.940 ;
        RECT  12.615 2.550 12.875 3.940 ;
        RECT  10.900 3.440 12.615 3.940 ;
        RECT  10.640 3.285 10.900 3.940 ;
        RECT  9.175 3.440 10.640 3.940 ;
        RECT  8.915 3.285 9.175 3.940 ;
        RECT  7.515 3.440 8.915 3.940 ;
        RECT  7.255 3.285 7.515 3.940 ;
        RECT  6.450 3.440 7.255 3.940 ;
        RECT  6.190 3.285 6.450 3.940 ;
        RECT  2.335 3.440 6.190 3.940 ;
        RECT  2.075 2.860 2.335 3.940 ;
        RECT  0.965 3.440 2.075 3.940 ;
        RECT  0.705 2.805 0.965 3.940 ;
        RECT  0.000 3.440 0.705 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.925 1.505 15.125 1.765 ;
        RECT  14.765 1.505 14.925 2.745 ;
        RECT  13.440 2.585 14.765 2.745 ;
        RECT  13.415 1.015 13.440 2.745 ;
        RECT  13.280 1.015 13.415 3.025 ;
        RECT  13.270 1.015 13.280 1.175 ;
        RECT  13.155 2.085 13.280 3.025 ;
        RECT  13.010 0.575 13.270 1.175 ;
        RECT  12.440 2.130 13.155 2.290 ;
        RECT  12.890 1.550 13.100 1.810 ;
        RECT  12.840 1.550 12.890 1.940 ;
        RECT  12.730 1.600 12.840 1.940 ;
        RECT  12.320 1.780 12.730 1.940 ;
        RECT  12.435 2.130 12.440 2.390 ;
        RECT  12.275 2.130 12.435 3.105 ;
        RECT  12.160 0.715 12.320 1.940 ;
        RECT  5.975 2.945 12.275 3.105 ;
        RECT  11.565 0.715 12.160 0.875 ;
        RECT  12.095 1.780 12.160 1.940 ;
        RECT  11.935 1.780 12.095 2.540 ;
        RECT  11.820 1.065 11.980 1.595 ;
        RECT  11.800 2.380 11.935 2.540 ;
        RECT  11.755 1.435 11.820 1.595 ;
        RECT  11.540 2.380 11.800 2.755 ;
        RECT  11.595 1.435 11.755 2.025 ;
        RECT  11.585 1.865 11.595 2.025 ;
        RECT  11.325 1.865 11.585 2.125 ;
        RECT  11.305 0.715 11.565 1.230 ;
        RECT  9.990 2.380 11.540 2.540 ;
        RECT  11.140 1.410 11.410 1.590 ;
        RECT  10.210 1.915 11.325 2.075 ;
        RECT  9.890 1.070 11.305 1.230 ;
        RECT  9.720 1.410 11.140 1.570 ;
        RECT  9.950 1.750 10.210 2.075 ;
        RECT  9.830 2.330 9.990 2.590 ;
        RECT  9.650 1.915 9.950 2.075 ;
        RECT  9.630 0.845 9.890 1.230 ;
        RECT  9.330 1.410 9.720 1.670 ;
        RECT  9.490 1.915 9.650 2.760 ;
        RECT  5.990 2.600 9.490 2.760 ;
        RECT  9.305 1.135 9.330 1.670 ;
        RECT  9.145 1.135 9.305 2.415 ;
        RECT  8.560 1.135 9.145 1.295 ;
        RECT  8.340 2.255 9.145 2.415 ;
        RECT  8.805 1.515 8.965 1.775 ;
        RECT  8.075 1.570 8.805 1.730 ;
        RECT  8.460 0.775 8.560 1.295 ;
        RECT  8.400 0.585 8.460 1.295 ;
        RECT  8.300 0.585 8.400 1.035 ;
        RECT  5.970 0.585 8.300 0.745 ;
        RECT  7.915 1.175 8.075 2.355 ;
        RECT  7.910 1.175 7.915 1.335 ;
        RECT  6.340 2.195 7.915 2.355 ;
        RECT  7.650 1.075 7.910 1.335 ;
        RECT  7.470 1.675 7.685 1.935 ;
        RECT  7.425 0.930 7.470 1.935 ;
        RECT  7.310 0.930 7.425 1.835 ;
        RECT  5.540 0.930 7.310 1.090 ;
        RECT  6.275 1.270 6.810 1.430 ;
        RECT  6.180 2.140 6.340 2.400 ;
        RECT  6.115 1.270 6.275 1.615 ;
        RECT  5.855 1.455 6.115 1.615 ;
        RECT  5.855 2.245 5.990 2.760 ;
        RECT  5.815 2.945 5.975 3.215 ;
        RECT  5.810 0.485 5.970 0.745 ;
        RECT  5.830 1.455 5.855 2.760 ;
        RECT  5.695 1.455 5.830 2.405 ;
        RECT  4.615 3.055 5.815 3.215 ;
        RECT  5.480 0.485 5.810 0.645 ;
        RECT  5.045 1.455 5.695 1.615 ;
        RECT  5.645 2.245 5.695 2.405 ;
        RECT  5.425 2.585 5.645 2.845 ;
        RECT  5.440 0.830 5.540 1.090 ;
        RECT  5.280 0.830 5.440 1.275 ;
        RECT  5.385 1.875 5.425 2.845 ;
        RECT  5.265 1.875 5.385 2.745 ;
        RECT  4.850 1.115 5.280 1.275 ;
        RECT  4.850 1.875 5.265 2.035 ;
        RECT  4.800 2.275 5.060 2.875 ;
        RECT  4.875 0.770 5.000 0.930 ;
        RECT  4.715 0.475 4.875 0.930 ;
        RECT  4.690 1.115 4.850 2.035 ;
        RECT  3.415 2.395 4.800 2.555 ;
        RECT  3.160 0.475 4.715 0.635 ;
        RECT  4.060 1.205 4.320 1.465 ;
        RECT  3.945 2.735 4.105 2.995 ;
        RECT  3.550 0.835 4.060 0.995 ;
        RECT  4.015 1.255 4.060 1.465 ;
        RECT  3.855 1.255 4.015 2.205 ;
        RECT  3.785 2.735 3.945 3.205 ;
        RECT  1.770 1.255 3.855 1.415 ;
        RECT  3.675 2.045 3.855 2.205 ;
        RECT  2.690 3.045 3.785 3.205 ;
        RECT  3.390 0.835 3.550 1.075 ;
        RECT  3.255 2.395 3.415 2.760 ;
        RECT  2.110 0.915 3.390 1.075 ;
        RECT  3.225 2.600 3.255 2.760 ;
        RECT  2.965 2.600 3.225 2.860 ;
        RECT  2.900 0.475 3.160 0.735 ;
        RECT  1.935 2.175 3.015 2.335 ;
        RECT  2.530 2.520 2.690 3.205 ;
        RECT  1.765 2.520 2.530 2.680 ;
        RECT  1.950 0.635 2.110 1.075 ;
        RECT  1.935 1.600 1.985 1.760 ;
        RECT  1.635 0.635 1.950 0.795 ;
        RECT  1.725 1.600 1.935 2.335 ;
        RECT  1.610 0.975 1.770 1.415 ;
        RECT  1.605 2.520 1.765 3.055 ;
        RECT  1.395 2.175 1.725 2.335 ;
        RECT  1.375 0.535 1.635 0.795 ;
        RECT  0.385 0.975 1.610 1.135 ;
        RECT  1.505 2.795 1.605 3.055 ;
        RECT  0.785 1.315 1.395 1.475 ;
        RECT  1.185 2.175 1.395 2.545 ;
        RECT  1.135 2.285 1.185 2.545 ;
        RECT  0.785 2.285 1.135 2.445 ;
        RECT  0.625 1.315 0.785 2.445 ;
        RECT  0.335 0.975 0.385 1.295 ;
        RECT  0.335 2.080 0.385 2.340 ;
        RECT  0.175 0.975 0.335 2.340 ;
        RECT  0.125 0.975 0.175 1.295 ;
        RECT  0.125 2.080 0.175 2.340 ;
    END
END SEDFFX4

MACRO SEDFFX2
    CLASS CORE ;
    FOREIGN SEDFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.800 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.655 2.635 1.990 ;
        RECT  2.270 1.655 2.425 1.985 ;
        RECT  2.200 1.655 2.270 1.880 ;
        END
        ANTENNAGATEAREA     0.0676 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.700 1.510 1.990 ;
        END
        ANTENNAGATEAREA     0.1222 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.465 0.590 13.675 3.030 ;
        RECT  13.415 0.590 13.465 1.190 ;
        RECT  13.415 2.090 13.465 3.030 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.655 1.700 12.755 2.175 ;
        RECT  12.560 1.700 12.655 2.335 ;
        RECT  12.560 0.490 12.610 0.750 ;
        RECT  12.400 0.490 12.560 2.335 ;
        RECT  12.350 0.490 12.400 0.750 ;
        RECT  12.395 1.765 12.400 2.335 ;
        END
        ANTENNADIFFAREA     0.5803 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.650 0.525 3.050 ;
        RECT  0.265 2.520 0.335 3.050 ;
        RECT  0.125 2.520 0.265 2.810 ;
        END
        ANTENNAGATEAREA     0.1222 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.245 1.610 3.470 1.865 ;
        RECT  3.080 1.610 3.245 1.990 ;
        RECT  2.885 1.700 3.080 1.990 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.400 1.675 6.890 1.990 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.165 -0.250 13.800 0.250 ;
        RECT  12.905 -0.250 13.165 1.190 ;
        RECT  11.800 -0.250 12.905 0.250 ;
        RECT  11.540 -0.250 11.800 0.405 ;
        RECT  10.540 -0.250 11.540 0.250 ;
        RECT  10.280 -0.250 10.540 0.405 ;
        RECT  8.725 -0.250 10.280 0.250 ;
        RECT  8.465 -0.250 8.725 0.405 ;
        RECT  7.200 -0.250 8.465 0.250 ;
        RECT  6.260 -0.250 7.200 0.655 ;
        RECT  2.520 -0.250 6.260 0.250 ;
        RECT  2.260 -0.250 2.520 0.735 ;
        RECT  0.965 -0.250 2.260 0.250 ;
        RECT  0.705 -0.250 0.965 0.710 ;
        RECT  0.000 -0.250 0.705 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.165 3.440 13.800 3.940 ;
        RECT  12.905 2.930 13.165 3.940 ;
        RECT  11.820 3.440 12.905 3.940 ;
        RECT  11.560 3.285 11.820 3.940 ;
        RECT  10.980 3.440 11.560 3.940 ;
        RECT  10.380 3.285 10.980 3.940 ;
        RECT  8.920 3.440 10.380 3.940 ;
        RECT  7.980 3.285 8.920 3.940 ;
        RECT  7.180 3.440 7.980 3.940 ;
        RECT  6.100 3.285 7.180 3.940 ;
        RECT  2.345 3.440 6.100 3.940 ;
        RECT  2.085 2.875 2.345 3.940 ;
        RECT  0.965 3.440 2.085 3.940 ;
        RECT  0.705 2.760 0.965 3.940 ;
        RECT  0.000 3.440 0.705 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.125 1.505 13.285 1.765 ;
        RECT  13.095 1.605 13.125 1.765 ;
        RECT  12.935 1.605 13.095 2.745 ;
        RECT  12.220 2.585 12.935 2.745 ;
        RECT  12.210 2.585 12.220 2.870 ;
        RECT  12.050 1.000 12.210 2.870 ;
        RECT  11.950 1.000 12.050 1.260 ;
        RECT  11.960 2.530 12.050 2.870 ;
        RECT  11.415 2.530 11.960 2.690 ;
        RECT  11.505 1.545 11.870 1.810 ;
        RECT  11.345 1.100 11.505 2.310 ;
        RECT  11.255 2.530 11.415 3.125 ;
        RECT  10.910 1.100 11.345 1.260 ;
        RECT  11.080 2.150 11.345 2.310 ;
        RECT  11.155 2.865 11.255 3.125 ;
        RECT  5.760 2.890 11.155 3.050 ;
        RECT  10.995 1.480 11.095 1.740 ;
        RECT  10.980 2.150 11.080 2.410 ;
        RECT  10.835 1.480 10.995 1.940 ;
        RECT  10.820 2.150 10.980 2.625 ;
        RECT  10.650 1.000 10.910 1.260 ;
        RECT  9.950 1.780 10.835 1.940 ;
        RECT  9.730 2.465 10.820 2.625 ;
        RECT  9.680 1.000 10.650 1.160 ;
        RECT  9.785 1.780 9.950 2.190 ;
        RECT  9.250 1.340 9.850 1.600 ;
        RECT  9.390 1.930 9.785 2.190 ;
        RECT  9.570 2.415 9.730 2.675 ;
        RECT  9.420 0.795 9.680 1.160 ;
        RECT  9.350 1.930 9.390 2.705 ;
        RECT  9.230 2.030 9.350 2.705 ;
        RECT  9.065 1.340 9.250 1.500 ;
        RECT  6.720 2.545 9.230 2.705 ;
        RECT  9.045 1.235 9.065 1.500 ;
        RECT  8.885 1.235 9.045 2.360 ;
        RECT  8.230 1.235 8.885 1.395 ;
        RECT  8.450 2.200 8.885 2.360 ;
        RECT  8.445 1.620 8.705 1.880 ;
        RECT  8.185 2.125 8.450 2.360 ;
        RECT  7.865 1.670 8.445 1.830 ;
        RECT  8.070 0.430 8.230 1.395 ;
        RECT  7.430 0.430 8.070 0.590 ;
        RECT  7.705 1.175 7.865 2.330 ;
        RECT  7.510 1.175 7.705 1.435 ;
        RECT  6.220 2.170 7.705 2.330 ;
        RECT  7.265 1.675 7.525 1.935 ;
        RECT  7.250 1.675 7.265 1.835 ;
        RECT  7.090 0.880 7.250 1.835 ;
        RECT  5.540 0.880 7.090 1.040 ;
        RECT  6.460 2.510 6.720 2.705 ;
        RECT  6.045 1.225 6.570 1.385 ;
        RECT  5.760 2.545 6.460 2.705 ;
        RECT  6.150 1.910 6.220 2.330 ;
        RECT  6.060 1.810 6.150 2.330 ;
        RECT  5.890 1.810 6.060 2.070 ;
        RECT  5.885 1.225 6.045 1.605 ;
        RECT  5.620 1.445 5.885 1.605 ;
        RECT  5.620 2.245 5.760 2.705 ;
        RECT  5.600 2.890 5.760 3.215 ;
        RECT  5.600 1.445 5.620 2.705 ;
        RECT  5.460 1.445 5.600 2.405 ;
        RECT  4.470 3.055 5.600 3.215 ;
        RECT  5.440 0.750 5.540 1.040 ;
        RECT  5.020 1.445 5.460 1.605 ;
        RECT  5.410 2.245 5.460 2.405 ;
        RECT  5.280 0.750 5.440 1.265 ;
        RECT  5.220 2.615 5.405 2.775 ;
        RECT  4.820 1.105 5.280 1.265 ;
        RECT  5.060 1.875 5.220 2.775 ;
        RECT  4.820 1.875 5.060 2.035 ;
        RECT  4.710 0.575 4.970 0.925 ;
        RECT  4.685 2.445 4.845 2.825 ;
        RECT  4.660 1.105 4.820 2.035 ;
        RECT  3.130 0.575 4.710 0.735 ;
        RECT  3.385 2.445 4.685 2.605 ;
        RECT  3.985 1.260 4.290 1.525 ;
        RECT  3.945 2.785 4.045 3.045 ;
        RECT  2.080 0.915 4.030 1.075 ;
        RECT  3.825 1.260 3.985 2.265 ;
        RECT  3.785 2.785 3.945 3.205 ;
        RECT  1.740 1.260 3.825 1.420 ;
        RECT  3.585 2.105 3.825 2.265 ;
        RECT  2.690 3.045 3.785 3.205 ;
        RECT  3.225 2.445 3.385 2.860 ;
        RECT  2.935 2.700 3.225 2.860 ;
        RECT  2.870 0.475 3.130 0.735 ;
        RECT  1.935 2.175 3.025 2.335 ;
        RECT  2.530 2.535 2.690 3.205 ;
        RECT  1.740 2.535 2.530 2.695 ;
        RECT  1.920 0.550 2.080 1.075 ;
        RECT  1.935 1.600 1.985 1.760 ;
        RECT  1.885 1.600 1.935 2.335 ;
        RECT  1.605 0.550 1.920 0.710 ;
        RECT  1.725 1.600 1.885 2.345 ;
        RECT  1.580 0.890 1.740 1.420 ;
        RECT  1.580 2.535 1.740 3.020 ;
        RECT  1.395 2.185 1.725 2.345 ;
        RECT  1.345 0.450 1.605 0.710 ;
        RECT  0.385 0.890 1.580 1.050 ;
        RECT  1.480 2.760 1.580 3.020 ;
        RECT  0.785 1.230 1.395 1.390 ;
        RECT  1.185 2.185 1.395 2.505 ;
        RECT  1.135 2.245 1.185 2.505 ;
        RECT  0.785 2.245 1.135 2.405 ;
        RECT  0.625 1.230 0.785 2.405 ;
        RECT  0.335 0.890 0.385 1.290 ;
        RECT  0.335 2.065 0.385 2.325 ;
        RECT  0.225 0.890 0.335 2.325 ;
        RECT  0.175 1.030 0.225 2.325 ;
        RECT  0.125 1.030 0.175 1.290 ;
        RECT  0.125 2.065 0.175 2.325 ;
    END
END SEDFFX2

MACRO SEDFFX1
    CLASS CORE ;
    FOREIGN SEDFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 1.610 2.265 1.990 ;
        END
        ANTENNAGATEAREA     0.0429 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.645 1.300 1.990 ;
        END
        ANTENNAGATEAREA     0.0949 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.375 0.575 11.395 2.745 ;
        RECT  11.235 0.575 11.375 2.810 ;
        RECT  11.115 0.575 11.235 0.835 ;
        RECT  11.165 2.135 11.235 2.810 ;
        RECT  11.115 2.135 11.165 2.735 ;
        END
        ANTENNADIFFAREA     0.4414 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.915 1.015 11.055 1.955 ;
        RECT  10.895 1.015 10.915 2.585 ;
        RECT  10.855 1.015 10.895 1.175 ;
        RECT  10.865 1.795 10.895 2.585 ;
        RECT  10.755 1.795 10.865 2.810 ;
        RECT  10.695 0.640 10.855 1.175 ;
        RECT  10.705 2.110 10.755 2.810 ;
        RECT  10.315 2.650 10.705 2.810 ;
        RECT  10.355 0.640 10.695 0.800 ;
        RECT  10.095 0.540 10.355 0.800 ;
        RECT  10.055 2.650 10.315 3.065 ;
        END
        ANTENNADIFFAREA     0.3332 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 2.520 0.795 2.810 ;
        RECT  0.255 2.550 0.585 2.810 ;
        END
        ANTENNAGATEAREA     0.0949 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.750 1.665 3.155 1.990 ;
        END
        ANTENNAGATEAREA     0.0455 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 2.110 6.775 2.400 ;
        RECT  6.565 1.875 6.725 2.400 ;
        RECT  6.150 1.875 6.565 2.035 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.865 -0.250 11.500 0.250 ;
        RECT  10.605 -0.250 10.865 0.405 ;
        RECT  9.795 -0.250 10.605 0.250 ;
        RECT  9.535 -0.250 9.795 0.405 ;
        RECT  8.245 -0.250 9.535 0.250 ;
        RECT  7.985 -0.250 8.245 1.015 ;
        RECT  6.555 -0.250 7.985 0.250 ;
        RECT  5.955 -0.250 6.555 0.590 ;
        RECT  2.365 -0.250 5.955 0.250 ;
        RECT  2.205 -0.250 2.365 0.705 ;
        RECT  0.965 -0.250 2.205 0.250 ;
        RECT  0.705 -0.250 0.965 0.405 ;
        RECT  0.000 -0.250 0.705 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.165 3.440 11.500 3.940 ;
        RECT  10.565 3.285 11.165 3.940 ;
        RECT  9.805 3.440 10.565 3.940 ;
        RECT  9.545 2.955 9.805 3.940 ;
        RECT  8.100 3.440 9.545 3.940 ;
        RECT  7.460 3.285 8.100 3.940 ;
        RECT  6.535 3.440 7.460 3.940 ;
        RECT  5.885 3.285 6.535 3.940 ;
        RECT  2.045 3.440 5.885 3.940 ;
        RECT  1.785 2.855 2.045 3.940 ;
        RECT  0.965 3.440 1.785 3.940 ;
        RECT  0.705 2.990 0.965 3.940 ;
        RECT  0.000 3.440 0.705 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.505 1.355 10.715 1.615 ;
        RECT  10.345 1.085 10.505 2.310 ;
        RECT  10.135 1.085 10.345 1.345 ;
        RECT  10.090 2.045 10.345 2.310 ;
        RECT  9.885 1.590 10.145 1.850 ;
        RECT  9.640 2.150 10.090 2.310 ;
        RECT  8.995 1.690 9.885 1.850 ;
        RECT  9.380 2.075 9.640 2.335 ;
        RECT  9.335 2.175 9.380 2.335 ;
        RECT  9.175 2.175 9.335 3.105 ;
        RECT  8.625 0.430 9.205 0.590 ;
        RECT  4.485 2.945 9.175 3.105 ;
        RECT  8.995 0.860 9.065 1.120 ;
        RECT  8.835 0.860 8.995 2.705 ;
        RECT  8.805 0.860 8.835 1.120 ;
        RECT  8.750 2.445 8.835 2.705 ;
        RECT  8.570 0.430 8.625 2.000 ;
        RECT  8.465 0.430 8.570 2.765 ;
        RECT  8.410 1.750 8.465 2.765 ;
        RECT  6.135 2.605 8.410 2.765 ;
        RECT  8.070 1.195 8.230 2.425 ;
        RECT  7.675 1.195 8.070 1.355 ;
        RECT  7.475 2.265 8.070 2.425 ;
        RECT  7.115 1.895 7.890 2.055 ;
        RECT  7.575 0.655 7.675 1.355 ;
        RECT  7.515 0.430 7.575 1.355 ;
        RECT  7.415 0.430 7.515 0.915 ;
        RECT  6.995 0.430 7.415 0.590 ;
        RECT  7.125 1.165 7.285 1.695 ;
        RECT  7.115 1.535 7.125 1.695 ;
        RECT  6.955 1.535 7.115 2.425 ;
        RECT  5.930 1.535 6.955 1.695 ;
        RECT  6.580 1.195 6.945 1.355 ;
        RECT  6.420 0.790 6.580 1.355 ;
        RECT  5.235 0.790 6.420 0.950 ;
        RECT  5.875 2.260 6.135 2.765 ;
        RECT  5.490 1.150 6.130 1.310 ;
        RECT  5.670 1.490 5.930 1.750 ;
        RECT  5.490 2.260 5.875 2.420 ;
        RECT  5.330 1.150 5.490 2.420 ;
        RECT  5.245 1.245 5.330 2.295 ;
        RECT  5.055 2.600 5.255 2.760 ;
        RECT  4.765 1.245 5.245 1.505 ;
        RECT  5.135 0.690 5.235 0.950 ;
        RECT  4.975 0.690 5.135 1.065 ;
        RECT  4.895 2.075 5.055 2.760 ;
        RECT  4.445 0.905 4.975 1.065 ;
        RECT  4.445 2.075 4.895 2.235 ;
        RECT  3.050 2.430 4.685 2.590 ;
        RECT  4.395 0.445 4.655 0.705 ;
        RECT  4.225 2.770 4.485 3.105 ;
        RECT  4.285 0.905 4.445 2.235 ;
        RECT  3.165 0.545 4.395 0.705 ;
        RECT  3.495 1.295 4.105 1.455 ;
        RECT  2.025 0.925 3.905 1.085 ;
        RECT  3.545 2.770 3.805 3.060 ;
        RECT  3.495 2.085 3.605 2.245 ;
        RECT  2.425 2.900 3.545 3.060 ;
        RECT  3.335 1.265 3.495 2.245 ;
        RECT  1.685 1.265 3.335 1.425 ;
        RECT  2.905 0.445 3.165 0.705 ;
        RECT  2.890 2.430 3.050 2.710 ;
        RECT  2.665 2.550 2.890 2.710 ;
        RECT  1.715 2.170 2.725 2.330 ;
        RECT  2.265 2.515 2.425 3.060 ;
        RECT  1.475 2.515 2.265 2.675 ;
        RECT  1.865 0.430 2.025 1.085 ;
        RECT  1.575 0.430 1.865 0.590 ;
        RECT  1.555 1.630 1.715 2.330 ;
        RECT  1.525 0.770 1.685 1.425 ;
        RECT  0.725 2.170 1.555 2.330 ;
        RECT  0.385 0.770 1.525 0.930 ;
        RECT  1.315 2.515 1.475 2.950 ;
        RECT  1.185 1.110 1.345 1.390 ;
        RECT  1.215 2.690 1.315 2.950 ;
        RECT  0.725 1.230 1.185 1.390 ;
        RECT  0.565 1.230 0.725 2.330 ;
        RECT  0.225 0.770 0.385 2.310 ;
        RECT  0.125 1.030 0.225 2.310 ;
    END
END SEDFFX1

MACRO SEDFFXL
    CLASS CORE ;
    FOREIGN SEDFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 1.610 2.265 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.645 1.300 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.215 0.650 11.375 2.810 ;
        RECT  11.115 0.650 11.215 0.910 ;
        RECT  11.165 2.210 11.215 2.810 ;
        RECT  11.115 2.210 11.165 2.470 ;
        END
        ANTENNADIFFAREA     0.2528 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.915 1.090 11.025 2.030 ;
        RECT  10.865 1.090 10.915 2.945 ;
        RECT  10.780 1.090 10.865 1.250 ;
        RECT  10.755 1.870 10.865 2.945 ;
        RECT  10.620 0.805 10.780 1.250 ;
        RECT  10.705 2.110 10.755 2.945 ;
        RECT  10.260 2.785 10.705 2.945 ;
        RECT  10.415 0.805 10.620 0.965 ;
        RECT  10.155 0.705 10.415 0.965 ;
        RECT  10.000 2.785 10.260 3.045 ;
        END
        ANTENNADIFFAREA     0.2320 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 2.520 0.795 2.810 ;
        RECT  0.255 2.550 0.585 2.810 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.750 1.615 3.155 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 2.110 6.775 2.400 ;
        RECT  6.485 2.110 6.565 2.335 ;
        RECT  6.325 1.875 6.485 2.335 ;
        RECT  6.225 1.875 6.325 2.035 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.850 -0.250 11.500 0.250 ;
        RECT  10.590 -0.250 10.850 0.405 ;
        RECT  9.785 -0.250 10.590 0.250 ;
        RECT  9.525 -0.250 9.785 0.405 ;
        RECT  8.195 -0.250 9.525 0.250 ;
        RECT  7.935 -0.250 8.195 1.015 ;
        RECT  6.555 -0.250 7.935 0.250 ;
        RECT  5.955 -0.250 6.555 0.590 ;
        RECT  2.365 -0.250 5.955 0.250 ;
        RECT  2.205 -0.250 2.365 0.705 ;
        RECT  0.965 -0.250 2.205 0.250 ;
        RECT  0.705 -0.250 0.965 0.405 ;
        RECT  0.000 -0.250 0.705 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.860 3.440 11.500 3.940 ;
        RECT  10.600 3.285 10.860 3.940 ;
        RECT  9.700 3.440 10.600 3.940 ;
        RECT  9.440 2.830 9.700 3.940 ;
        RECT  8.095 3.440 9.440 3.940 ;
        RECT  7.465 3.285 8.095 3.940 ;
        RECT  6.585 3.440 7.465 3.940 ;
        RECT  5.885 3.285 6.585 3.940 ;
        RECT  2.045 3.440 5.885 3.940 ;
        RECT  1.785 2.855 2.045 3.940 ;
        RECT  0.965 3.440 1.785 3.940 ;
        RECT  0.705 2.990 0.965 3.940 ;
        RECT  0.000 3.440 0.705 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.380 1.430 10.685 1.690 ;
        RECT  10.290 1.215 10.380 2.290 ;
        RECT  10.220 1.215 10.290 2.470 ;
        RECT  10.105 1.215 10.220 1.475 ;
        RECT  10.030 2.130 10.220 2.470 ;
        RECT  9.880 1.690 10.040 1.950 ;
        RECT  9.470 2.130 10.030 2.290 ;
        RECT  9.720 0.865 9.880 1.925 ;
        RECT  9.045 0.865 9.720 1.025 ;
        RECT  9.250 1.605 9.470 2.290 ;
        RECT  9.210 1.605 9.250 3.105 ;
        RECT  9.090 2.130 9.210 3.105 ;
        RECT  8.570 0.525 9.205 0.685 ;
        RECT  4.485 2.945 9.090 3.105 ;
        RECT  8.910 0.865 9.045 1.125 ;
        RECT  8.750 0.865 8.910 2.765 ;
        RECT  8.525 0.525 8.570 1.480 ;
        RECT  8.410 0.525 8.525 2.765 ;
        RECT  8.365 1.320 8.410 2.765 ;
        RECT  6.135 2.605 8.365 2.765 ;
        RECT  8.025 1.195 8.185 2.425 ;
        RECT  7.625 1.195 8.025 1.355 ;
        RECT  7.475 2.265 8.025 2.425 ;
        RECT  7.115 1.895 7.845 2.055 ;
        RECT  7.465 0.430 7.625 1.355 ;
        RECT  6.995 0.430 7.465 0.690 ;
        RECT  7.125 1.160 7.285 1.695 ;
        RECT  7.115 1.535 7.125 1.695 ;
        RECT  6.955 1.535 7.115 2.405 ;
        RECT  5.880 1.535 6.955 1.695 ;
        RECT  6.580 1.195 6.945 1.355 ;
        RECT  6.420 0.810 6.580 1.355 ;
        RECT  5.020 0.810 6.420 0.970 ;
        RECT  6.045 2.215 6.135 2.765 ;
        RECT  5.405 1.155 6.130 1.315 ;
        RECT  5.875 2.135 6.045 2.765 ;
        RECT  5.720 1.535 5.880 1.865 ;
        RECT  5.405 2.135 5.875 2.295 ;
        RECT  5.245 1.155 5.405 2.295 ;
        RECT  5.055 2.500 5.255 2.760 ;
        RECT  4.765 1.245 5.245 1.505 ;
        RECT  4.895 1.685 5.055 2.760 ;
        RECT  4.860 0.810 5.020 0.995 ;
        RECT  4.445 1.685 4.895 1.845 ;
        RECT  4.445 0.835 4.860 0.995 ;
        RECT  4.425 2.330 4.685 2.590 ;
        RECT  2.905 0.495 4.645 0.655 ;
        RECT  4.225 2.770 4.485 3.105 ;
        RECT  4.285 0.835 4.445 1.845 ;
        RECT  3.050 2.430 4.425 2.590 ;
        RECT  3.495 1.295 4.105 1.455 ;
        RECT  2.025 0.925 3.905 1.085 ;
        RECT  3.545 2.770 3.805 3.085 ;
        RECT  3.495 2.085 3.605 2.245 ;
        RECT  2.425 2.925 3.545 3.085 ;
        RECT  3.335 1.265 3.495 2.245 ;
        RECT  1.685 1.265 3.335 1.425 ;
        RECT  2.890 2.430 3.050 2.735 ;
        RECT  2.665 2.575 2.890 2.735 ;
        RECT  1.715 2.170 2.725 2.330 ;
        RECT  2.265 2.515 2.425 3.085 ;
        RECT  1.475 2.515 2.265 2.675 ;
        RECT  1.865 0.430 2.025 1.085 ;
        RECT  1.575 0.430 1.865 0.590 ;
        RECT  1.555 1.630 1.715 2.330 ;
        RECT  1.525 0.770 1.685 1.425 ;
        RECT  0.725 2.170 1.555 2.330 ;
        RECT  0.385 0.770 1.525 0.930 ;
        RECT  1.315 2.515 1.475 2.950 ;
        RECT  1.185 1.110 1.345 1.390 ;
        RECT  1.215 2.690 1.315 2.950 ;
        RECT  0.725 1.230 1.185 1.390 ;
        RECT  0.565 1.230 0.725 2.330 ;
        RECT  0.225 0.770 0.385 2.310 ;
        RECT  0.125 1.030 0.225 1.290 ;
        RECT  0.125 2.050 0.225 2.310 ;
    END
END SEDFFXL

MACRO SDFFTRX4
    CLASS CORE ;
    FOREIGN SDFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.340 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.700 4.015 2.015 ;
        RECT  3.420 1.755 3.805 2.015 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.375 1.725 2.535 2.340 ;
        RECT  1.275 2.180 2.375 2.340 ;
        RECT  1.115 1.850 1.275 2.340 ;
        RECT  0.795 1.850 1.115 2.010 ;
        RECT  0.775 1.515 0.795 2.010 ;
        RECT  0.585 1.460 0.775 2.010 ;
        RECT  0.505 1.460 0.585 1.720 ;
        END
        ANTENNAGATEAREA     0.3640 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.600 1.285 3.940 1.445 ;
        RECT  3.440 0.585 3.600 1.445 ;
        RECT  3.005 0.585 3.440 0.745 ;
        RECT  2.845 0.470 3.005 0.745 ;
        RECT  1.530 0.470 2.845 0.630 ;
        RECT  1.385 0.470 1.530 0.760 ;
        RECT  1.255 0.470 1.385 1.415 ;
        RECT  1.225 0.470 1.255 1.580 ;
        RECT  1.145 1.255 1.225 1.580 ;
        RECT  0.985 1.255 1.145 1.670 ;
        END
        ANTENNAGATEAREA     0.2028 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.410 0.570 11.670 2.215 ;
        RECT  11.165 1.290 11.410 1.990 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.205 1.290 13.215 2.175 ;
        RECT  13.005 1.015 13.205 2.305 ;
        RECT  12.690 1.015 13.005 1.215 ;
        RECT  12.755 2.105 13.005 2.305 ;
        RECT  12.690 2.105 12.755 2.585 ;
        RECT  12.430 0.595 12.690 1.215 ;
        RECT  12.430 2.105 12.690 3.045 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 1.595 1.940 1.990 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.650 1.290 4.935 1.735 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.200 -0.250 13.340 0.250 ;
        RECT  12.940 -0.250 13.200 0.795 ;
        RECT  12.180 -0.250 12.940 0.250 ;
        RECT  11.920 -0.250 12.180 1.270 ;
        RECT  11.120 -0.250 11.920 0.250 ;
        RECT  10.860 -0.250 11.120 0.405 ;
        RECT  10.170 -0.250 10.860 0.250 ;
        RECT  9.910 -0.250 10.170 0.855 ;
        RECT  8.370 -0.250 9.910 0.250 ;
        RECT  8.110 -0.250 8.370 0.405 ;
        RECT  7.310 -0.250 8.110 0.250 ;
        RECT  7.050 -0.250 7.310 0.405 ;
        RECT  4.495 -0.250 7.050 0.250 ;
        RECT  4.235 -0.250 4.495 0.405 ;
        RECT  3.585 -0.250 4.235 0.250 ;
        RECT  3.325 -0.250 3.585 0.405 ;
        RECT  1.025 -0.250 3.325 0.250 ;
        RECT  0.765 -0.250 1.025 1.075 ;
        RECT  0.000 -0.250 0.765 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.200 3.440 13.340 3.940 ;
        RECT  12.940 2.590 13.200 3.940 ;
        RECT  12.180 3.440 12.940 3.940 ;
        RECT  11.920 2.935 12.180 3.940 ;
        RECT  11.130 3.440 11.920 3.940 ;
        RECT  10.870 3.285 11.130 3.940 ;
        RECT  10.170 3.440 10.870 3.940 ;
        RECT  9.910 2.865 10.170 3.940 ;
        RECT  8.370 3.440 9.910 3.940 ;
        RECT  8.110 2.800 8.370 3.940 ;
        RECT  6.870 3.440 8.110 3.940 ;
        RECT  6.710 2.735 6.870 3.940 ;
        RECT  5.070 3.440 6.710 3.940 ;
        RECT  4.810 2.515 5.070 3.940 ;
        RECT  3.670 3.440 4.810 3.940 ;
        RECT  3.410 2.625 3.670 3.940 ;
        RECT  1.505 3.440 3.410 3.940 ;
        RECT  1.245 2.955 1.505 3.940 ;
        RECT  0.000 3.440 1.245 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.220 1.510 12.820 1.770 ;
        RECT  12.010 1.610 12.220 1.770 ;
        RECT  11.850 1.610 12.010 2.555 ;
        RECT  10.925 2.395 11.850 2.555 ;
        RECT  10.765 1.040 10.925 2.555 ;
        RECT  10.755 1.040 10.765 1.200 ;
        RECT  10.755 2.275 10.765 2.555 ;
        RECT  10.495 0.940 10.755 1.200 ;
        RECT  10.495 2.275 10.755 2.885 ;
        RECT  10.325 1.380 10.585 1.695 ;
        RECT  10.105 2.275 10.495 2.435 ;
        RECT  9.425 1.380 10.325 1.540 ;
        RECT  9.945 1.725 10.105 2.435 ;
        RECT  9.845 1.725 9.945 1.985 ;
        RECT  9.425 0.430 9.685 0.745 ;
        RECT  6.870 0.585 9.425 0.745 ;
        RECT  9.265 1.090 9.425 2.675 ;
        RECT  9.165 1.090 9.265 1.350 ;
        RECT  9.165 2.075 9.265 2.675 ;
        RECT  7.290 2.460 9.165 2.620 ;
        RECT  8.750 0.930 8.910 2.280 ;
        RECT  7.100 0.930 8.750 1.090 ;
        RECT  7.570 2.120 8.750 2.280 ;
        RECT  7.930 1.395 8.530 1.655 ;
        RECT  6.530 1.445 7.930 1.605 ;
        RECT  7.130 1.800 7.290 2.620 ;
        RECT  7.030 1.800 7.130 2.060 ;
        RECT  6.840 0.930 7.100 1.255 ;
        RECT  6.710 0.470 6.870 0.745 ;
        RECT  6.620 0.470 6.710 0.630 ;
        RECT  6.360 0.430 6.620 0.630 ;
        RECT  6.370 0.915 6.530 2.780 ;
        RECT  6.360 0.915 6.370 1.075 ;
        RECT  6.095 2.615 6.370 2.780 ;
        RECT  5.460 0.470 6.360 0.630 ;
        RECT  6.100 0.815 6.360 1.075 ;
        RECT  6.030 1.315 6.190 2.335 ;
        RECT  5.835 2.515 6.095 3.115 ;
        RECT  5.800 1.315 6.030 1.475 ;
        RECT  5.585 2.175 6.030 2.335 ;
        RECT  5.510 1.680 5.835 1.945 ;
        RECT  5.640 0.815 5.800 1.475 ;
        RECT  5.325 2.175 5.585 3.060 ;
        RECT  5.460 1.680 5.510 1.995 ;
        RECT  5.300 0.470 5.460 1.995 ;
        RECT  4.490 2.175 5.325 2.335 ;
        RECT  4.825 0.470 5.300 0.630 ;
        RECT  5.250 1.735 5.300 1.995 ;
        RECT  4.960 0.830 5.120 1.105 ;
        RECT  4.470 0.945 4.960 1.105 ;
        RECT  4.280 2.175 4.490 3.075 ;
        RECT  4.310 0.945 4.470 1.995 ;
        RECT  4.095 0.945 4.310 1.105 ;
        RECT  4.230 2.195 4.280 3.075 ;
        RECT  3.215 2.195 4.230 2.355 ;
        RECT  3.835 0.815 4.095 1.105 ;
        RECT  3.055 0.925 3.215 3.215 ;
        RECT  2.665 0.925 3.055 1.085 ;
        RECT  2.325 3.055 3.055 3.215 ;
        RECT  2.715 1.345 2.875 2.685 ;
        RECT  2.585 1.345 2.715 1.505 ;
        RECT  2.590 2.525 2.715 2.685 ;
        RECT  2.065 0.810 2.665 1.085 ;
        RECT  2.330 2.525 2.590 2.775 ;
        RECT  2.325 1.265 2.585 1.505 ;
        RECT  0.810 2.525 2.330 2.685 ;
        RECT  2.065 2.955 2.325 3.215 ;
        RECT  0.650 2.190 0.810 2.685 ;
        RECT  0.325 2.190 0.650 2.450 ;
        RECT  0.325 1.035 0.385 1.295 ;
        RECT  0.165 1.035 0.325 2.450 ;
        RECT  0.125 1.035 0.165 1.295 ;
    END
END SDFFTRX4

MACRO SDFFTRX2
    CLASS CORE ;
    FOREIGN SDFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.420 1.280 2.690 1.745 ;
        END
        ANTENNAGATEAREA     0.0806 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.530 1.490 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.2236 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.290 3.165 1.745 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.470 1.515 9.535 1.990 ;
        RECT  9.315 0.595 9.470 2.115 ;
        RECT  9.310 0.595 9.315 2.215 ;
        RECT  9.050 0.495 9.310 0.755 ;
        RECT  9.155 1.955 9.310 2.215 ;
        END
        ANTENNADIFFAREA     0.6779 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.195 0.600 10.455 3.045 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.995 1.475 1.255 1.990 ;
        END
        ANTENNAGATEAREA     0.1586 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.855 1.290 4.015 1.770 ;
        RECT  3.685 1.290 3.855 1.595 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.910 -0.250 10.580 0.250 ;
        RECT  9.650 -0.250 9.910 1.135 ;
        RECT  8.370 -0.250 9.650 0.250 ;
        RECT  8.110 -0.250 8.370 0.855 ;
        RECT  6.570 -0.250 8.110 0.250 ;
        RECT  6.310 -0.250 6.570 0.405 ;
        RECT  4.080 -0.250 6.310 0.250 ;
        RECT  3.820 -0.250 4.080 0.770 ;
        RECT  2.885 -0.250 3.820 0.250 ;
        RECT  2.625 -0.250 2.885 1.065 ;
        RECT  0.815 -0.250 2.625 0.250 ;
        RECT  0.555 -0.250 0.815 0.820 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.910 3.440 10.580 3.940 ;
        RECT  9.650 2.870 9.910 3.940 ;
        RECT  8.170 3.440 9.650 3.940 ;
        RECT  7.910 2.865 8.170 3.940 ;
        RECT  6.130 3.440 7.910 3.940 ;
        RECT  5.870 2.095 6.130 3.940 ;
        RECT  4.185 3.440 5.870 3.940 ;
        RECT  3.925 2.465 4.185 3.940 ;
        RECT  2.805 3.440 3.925 3.940 ;
        RECT  2.545 2.315 2.805 3.940 ;
        RECT  1.040 3.440 2.545 3.940 ;
        RECT  0.780 2.510 1.040 3.940 ;
        RECT  0.000 3.440 0.780 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.855 1.585 10.015 2.595 ;
        RECT  8.965 2.435 9.855 2.595 ;
        RECT  8.845 1.035 8.965 2.595 ;
        RECT  8.805 1.035 8.845 2.695 ;
        RECT  8.690 1.035 8.805 1.295 ;
        RECT  8.585 2.435 8.805 2.695 ;
        RECT  8.510 1.565 8.625 1.825 ;
        RECT  8.085 2.435 8.585 2.595 ;
        RECT  8.350 1.315 8.510 1.825 ;
        RECT  7.630 1.315 8.350 1.475 ;
        RECT  7.925 1.725 8.085 2.595 ;
        RECT  7.825 1.725 7.925 1.985 ;
        RECT  7.585 0.930 7.630 1.475 ;
        RECT  7.420 0.930 7.585 2.395 ;
        RECT  7.370 0.930 7.420 1.190 ;
        RECT  7.220 2.235 7.420 2.395 ;
        RECT  7.255 0.450 7.355 0.610 ;
        RECT  7.095 0.450 7.255 0.750 ;
        RECT  6.960 2.235 7.220 2.835 ;
        RECT  7.020 0.930 7.120 1.190 ;
        RECT  6.035 0.590 7.095 0.750 ;
        RECT  6.860 0.930 7.020 1.285 ;
        RECT  6.640 1.125 6.860 1.285 ;
        RECT  6.480 1.125 6.640 2.695 ;
        RECT  6.090 1.125 6.480 1.385 ;
        RECT  6.380 2.095 6.480 2.695 ;
        RECT  6.040 1.605 6.300 1.865 ;
        RECT  5.690 1.705 6.040 1.865 ;
        RECT  5.875 0.505 6.035 0.750 ;
        RECT  5.870 0.505 5.875 0.665 ;
        RECT  5.610 0.430 5.870 0.665 ;
        RECT  5.685 1.705 5.690 2.625 ;
        RECT  5.525 0.845 5.685 2.625 ;
        RECT  4.695 0.505 5.610 0.665 ;
        RECT  5.410 0.845 5.525 1.005 ;
        RECT  5.250 2.465 5.525 2.625 ;
        RECT  5.185 1.305 5.345 2.285 ;
        RECT  4.990 2.465 5.250 2.725 ;
        RECT  5.165 1.305 5.185 1.465 ;
        RECT  4.710 2.125 5.185 2.285 ;
        RECT  5.005 0.845 5.165 1.465 ;
        RECT  4.900 0.845 5.005 1.005 ;
        RECT  4.695 1.675 5.005 1.935 ;
        RECT  4.450 2.125 4.710 2.655 ;
        RECT  4.535 0.505 4.695 1.935 ;
        RECT  4.390 0.610 4.535 0.770 ;
        RECT  4.425 1.775 4.535 1.935 ;
        RECT  3.625 2.125 4.450 2.285 ;
        RECT  4.195 0.950 4.355 1.480 ;
        RECT  3.510 0.950 4.195 1.110 ;
        RECT  3.505 1.775 3.675 1.935 ;
        RECT  3.365 2.125 3.625 2.505 ;
        RECT  3.505 0.560 3.510 1.110 ;
        RECT  3.345 0.560 3.505 1.935 ;
        RECT  3.145 2.125 3.365 2.285 ;
        RECT  3.250 0.560 3.345 0.820 ;
        RECT  2.985 1.975 3.145 2.285 ;
        RECT  2.145 1.975 2.985 2.135 ;
        RECT  1.985 0.885 2.145 2.135 ;
        RECT  1.855 2.880 2.115 3.140 ;
        RECT  1.975 0.885 1.985 1.045 ;
        RECT  1.935 1.975 1.985 2.135 ;
        RECT  1.715 0.785 1.975 1.045 ;
        RECT  1.775 1.975 1.935 2.500 ;
        RECT  1.595 2.880 1.855 3.040 ;
        RECT  1.595 1.235 1.805 1.495 ;
        RECT  1.435 1.235 1.595 3.040 ;
        RECT  0.385 2.170 1.435 2.330 ;
        RECT  0.285 1.035 0.385 1.295 ;
        RECT  0.285 2.120 0.385 2.330 ;
        RECT  0.125 1.035 0.285 2.330 ;
    END
END SDFFTRX2

MACRO SDFFTRX1
    CLASS CORE ;
    FOREIGN SDFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 2.860 2.405 3.220 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 1.700 0.795 1.990 ;
        RECT  0.495 1.550 0.760 1.990 ;
        END
        ANTENNAGATEAREA     0.1456 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.110 1.300 3.165 1.560 ;
        RECT  2.740 1.290 3.110 1.585 ;
        END
        ANTENNAGATEAREA     0.0637 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.485 1.105 9.535 2.585 ;
        RECT  9.325 0.750 9.485 2.730 ;
        RECT  8.880 0.750 9.325 0.910 ;
        RECT  9.050 2.570 9.325 2.730 ;
        RECT  8.790 2.570 9.050 3.170 ;
        RECT  8.620 0.650 8.880 0.910 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.735 0.995 9.995 2.765 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.165 1.475 1.325 3.220 ;
        RECT  1.065 1.475 1.165 1.765 ;
        RECT  1.045 2.930 1.165 3.220 ;
        END
        ANTENNAGATEAREA     0.0832 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.855 1.290 4.015 1.770 ;
        RECT  3.685 1.290 3.855 1.600 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.435 -0.250 10.120 0.250 ;
        RECT  9.175 -0.250 9.435 0.405 ;
        RECT  8.270 -0.250 9.175 0.250 ;
        RECT  8.010 -0.250 8.270 0.855 ;
        RECT  6.620 -0.250 8.010 0.250 ;
        RECT  6.360 -0.250 6.620 0.405 ;
        RECT  4.080 -0.250 6.360 0.250 ;
        RECT  3.820 -0.250 4.080 0.770 ;
        RECT  2.885 -0.250 3.820 0.250 ;
        RECT  2.625 -0.250 2.885 0.975 ;
        RECT  0.815 -0.250 2.625 0.250 ;
        RECT  0.555 -0.250 0.815 0.820 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.600 3.440 10.120 3.940 ;
        RECT  9.340 3.285 9.600 3.940 ;
        RECT  7.960 3.440 9.340 3.940 ;
        RECT  7.700 2.845 7.960 3.940 ;
        RECT  6.160 3.440 7.700 3.940 ;
        RECT  5.900 2.255 6.160 3.940 ;
        RECT  4.185 3.440 5.900 3.940 ;
        RECT  3.925 2.515 4.185 3.940 ;
        RECT  2.745 3.440 3.925 3.940 ;
        RECT  2.585 2.245 2.745 3.940 ;
        RECT  0.855 3.440 2.585 3.940 ;
        RECT  0.855 2.180 0.955 2.440 ;
        RECT  0.695 2.180 0.855 3.940 ;
        RECT  0.000 3.440 0.695 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.990 1.880 9.145 2.140 ;
        RECT  8.830 1.320 8.990 2.385 ;
        RECT  8.800 1.320 8.830 1.480 ;
        RECT  8.540 2.225 8.830 2.385 ;
        RECT  8.640 1.195 8.800 1.480 ;
        RECT  8.460 1.785 8.650 2.045 ;
        RECT  8.280 2.225 8.540 2.820 ;
        RECT  8.300 1.315 8.460 2.045 ;
        RECT  7.525 1.315 8.300 1.475 ;
        RECT  8.120 2.225 8.280 2.385 ;
        RECT  7.960 1.870 8.120 2.385 ;
        RECT  7.365 1.035 7.525 2.565 ;
        RECT  7.265 1.035 7.365 1.295 ;
        RECT  7.220 2.405 7.365 2.565 ;
        RECT  6.160 0.690 7.355 0.850 ;
        RECT  6.960 2.405 7.220 2.665 ;
        RECT  6.915 1.030 7.015 1.290 ;
        RECT  6.755 1.030 6.915 1.595 ;
        RECT  6.670 1.435 6.755 1.595 ;
        RECT  6.670 2.485 6.710 2.745 ;
        RECT  6.510 1.435 6.670 2.745 ;
        RECT  6.240 1.435 6.510 1.595 ;
        RECT  6.450 2.485 6.510 2.745 ;
        RECT  6.070 1.815 6.330 2.075 ;
        RECT  5.980 1.335 6.240 1.595 ;
        RECT  6.000 0.475 6.160 0.850 ;
        RECT  5.685 1.915 6.070 2.075 ;
        RECT  5.880 0.475 6.000 0.635 ;
        RECT  5.670 0.470 5.880 0.635 ;
        RECT  5.685 0.845 5.730 1.005 ;
        RECT  5.525 0.845 5.685 2.675 ;
        RECT  4.720 0.470 5.670 0.630 ;
        RECT  5.470 0.845 5.525 1.005 ;
        RECT  5.280 2.515 5.525 2.675 ;
        RECT  5.290 1.305 5.345 2.335 ;
        RECT  5.185 0.810 5.290 2.335 ;
        RECT  5.020 2.515 5.280 2.775 ;
        RECT  5.130 0.810 5.185 1.465 ;
        RECT  4.710 2.175 5.185 2.335 ;
        RECT  4.900 0.810 5.130 1.060 ;
        RECT  4.720 1.685 5.005 1.945 ;
        RECT  4.685 0.470 4.720 1.945 ;
        RECT  4.450 2.175 4.710 2.655 ;
        RECT  4.560 0.470 4.685 1.995 ;
        RECT  4.390 0.610 4.560 0.770 ;
        RECT  4.425 1.735 4.560 1.995 ;
        RECT  3.675 2.175 4.450 2.335 ;
        RECT  4.195 0.950 4.355 1.480 ;
        RECT  3.510 0.950 4.195 1.110 ;
        RECT  3.505 1.785 3.675 1.945 ;
        RECT  3.415 2.175 3.675 2.505 ;
        RECT  3.505 0.560 3.510 1.110 ;
        RECT  3.345 0.560 3.505 1.945 ;
        RECT  3.105 2.175 3.415 2.335 ;
        RECT  3.250 0.560 3.345 0.820 ;
        RECT  2.945 1.885 3.105 2.335 ;
        RECT  2.405 1.885 2.945 2.045 ;
        RECT  2.245 0.795 2.405 2.475 ;
        RECT  2.005 0.795 2.245 0.955 ;
        RECT  1.915 2.315 2.245 2.475 ;
        RECT  1.905 1.135 2.065 2.135 ;
        RECT  1.745 0.695 2.005 0.955 ;
        RECT  1.655 2.315 1.915 2.575 ;
        RECT  0.385 1.135 1.905 1.295 ;
        RECT  0.285 1.035 0.385 1.295 ;
        RECT  0.285 2.180 0.385 2.440 ;
        RECT  0.125 1.035 0.285 2.440 ;
    END
END SDFFTRX1

MACRO SDFFTRXL
    CLASS CORE ;
    FOREIGN SDFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 2.860 2.405 3.220 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 1.700 0.795 1.990 ;
        RECT  0.495 1.550 0.760 1.990 ;
        END
        ANTENNAGATEAREA     0.1352 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.110 1.300 3.165 1.560 ;
        RECT  2.740 1.290 3.110 1.585 ;
        END
        ANTENNAGATEAREA     0.0559 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.485 1.105 9.535 2.585 ;
        RECT  9.325 0.750 9.485 2.900 ;
        RECT  8.935 0.750 9.325 0.910 ;
        RECT  9.045 2.740 9.325 2.900 ;
        RECT  8.785 2.740 9.045 3.000 ;
        RECT  8.675 0.650 8.935 0.910 ;
        END
        ANTENNADIFFAREA     0.2142 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.735 1.030 9.995 2.595 ;
        END
        ANTENNADIFFAREA     0.2142 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.165 1.475 1.325 3.225 ;
        RECT  1.065 1.475 1.165 1.765 ;
        RECT  1.070 2.930 1.165 3.225 ;
        RECT  1.045 2.930 1.070 3.220 ;
        END
        ANTENNAGATEAREA     0.0650 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.855 1.290 4.015 1.770 ;
        RECT  3.685 1.290 3.855 1.600 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.525 -0.250 10.120 0.250 ;
        RECT  9.265 -0.250 9.525 0.405 ;
        RECT  8.355 -0.250 9.265 0.250 ;
        RECT  8.095 -0.250 8.355 0.855 ;
        RECT  6.620 -0.250 8.095 0.250 ;
        RECT  6.360 -0.250 6.620 0.405 ;
        RECT  4.080 -0.250 6.360 0.250 ;
        RECT  3.820 -0.250 4.080 0.770 ;
        RECT  2.885 -0.250 3.820 0.250 ;
        RECT  2.625 -0.250 2.885 0.975 ;
        RECT  0.815 -0.250 2.625 0.250 ;
        RECT  0.555 -0.250 0.815 0.820 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.595 3.440 10.120 3.940 ;
        RECT  9.335 3.285 9.595 3.940 ;
        RECT  7.960 3.440 9.335 3.940 ;
        RECT  7.700 2.925 7.960 3.940 ;
        RECT  6.160 3.440 7.700 3.940 ;
        RECT  5.900 2.340 6.160 3.940 ;
        RECT  4.185 3.440 5.900 3.940 ;
        RECT  3.925 2.515 4.185 3.940 ;
        RECT  2.745 3.440 3.925 3.940 ;
        RECT  2.585 2.245 2.745 3.940 ;
        RECT  0.855 3.440 2.585 3.940 ;
        RECT  0.855 2.180 0.955 2.440 ;
        RECT  0.695 2.180 0.855 3.940 ;
        RECT  0.000 3.440 0.695 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.990 1.880 9.145 2.140 ;
        RECT  8.830 1.180 8.990 2.560 ;
        RECT  8.675 1.180 8.830 1.440 ;
        RECT  8.535 2.400 8.830 2.560 ;
        RECT  8.460 1.620 8.650 2.220 ;
        RECT  8.275 2.400 8.535 2.820 ;
        RECT  8.390 1.315 8.460 2.220 ;
        RECT  8.300 1.315 8.390 2.045 ;
        RECT  7.615 1.315 8.300 1.475 ;
        RECT  8.075 2.400 8.275 2.560 ;
        RECT  7.915 1.870 8.075 2.560 ;
        RECT  7.815 1.870 7.915 2.130 ;
        RECT  7.455 1.030 7.615 2.500 ;
        RECT  7.355 1.030 7.455 1.290 ;
        RECT  7.210 2.340 7.455 2.500 ;
        RECT  7.155 0.585 7.415 0.845 ;
        RECT  6.950 2.340 7.210 2.600 ;
        RECT  6.160 0.585 7.155 0.745 ;
        RECT  6.945 1.030 7.045 1.290 ;
        RECT  6.785 1.030 6.945 1.495 ;
        RECT  6.670 1.335 6.785 1.495 ;
        RECT  6.510 1.335 6.670 2.600 ;
        RECT  6.240 1.335 6.510 1.495 ;
        RECT  6.460 2.340 6.510 2.600 ;
        RECT  6.070 1.900 6.330 2.160 ;
        RECT  5.980 1.335 6.240 1.595 ;
        RECT  6.000 0.475 6.160 0.745 ;
        RECT  5.720 2.000 6.070 2.160 ;
        RECT  4.700 0.475 6.000 0.635 ;
        RECT  5.720 0.865 5.730 1.025 ;
        RECT  5.560 0.865 5.720 2.675 ;
        RECT  5.470 0.865 5.560 1.025 ;
        RECT  5.280 2.515 5.560 2.675 ;
        RECT  5.290 1.305 5.380 2.335 ;
        RECT  5.220 0.815 5.290 2.335 ;
        RECT  5.020 2.515 5.280 2.775 ;
        RECT  5.130 0.815 5.220 1.465 ;
        RECT  4.710 2.175 5.220 2.335 ;
        RECT  4.900 0.815 5.130 1.075 ;
        RECT  4.700 1.685 5.005 1.945 ;
        RECT  4.450 2.175 4.710 2.655 ;
        RECT  4.685 0.475 4.700 1.945 ;
        RECT  4.540 0.475 4.685 1.995 ;
        RECT  4.390 0.610 4.540 0.770 ;
        RECT  4.425 1.735 4.540 1.995 ;
        RECT  3.675 2.175 4.450 2.335 ;
        RECT  4.195 0.950 4.355 1.480 ;
        RECT  3.510 0.950 4.195 1.110 ;
        RECT  3.505 1.785 3.675 1.945 ;
        RECT  3.415 2.175 3.675 2.505 ;
        RECT  3.505 0.560 3.510 1.110 ;
        RECT  3.345 0.560 3.505 1.945 ;
        RECT  3.105 2.175 3.415 2.335 ;
        RECT  3.250 0.560 3.345 0.820 ;
        RECT  2.945 1.885 3.105 2.335 ;
        RECT  2.405 1.885 2.945 2.045 ;
        RECT  2.245 0.795 2.405 2.475 ;
        RECT  2.005 0.795 2.245 0.955 ;
        RECT  1.915 2.315 2.245 2.475 ;
        RECT  1.905 1.135 2.065 2.135 ;
        RECT  1.745 0.695 2.005 0.955 ;
        RECT  1.655 2.315 1.915 2.575 ;
        RECT  0.385 1.135 1.905 1.295 ;
        RECT  0.285 1.035 0.385 1.295 ;
        RECT  0.285 2.180 0.385 2.440 ;
        RECT  0.125 1.035 0.285 2.440 ;
    END
END SDFFTRXL

MACRO SDFFNSRX4
    CLASS CORE ;
    FOREIGN SDFFNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.975 2.930 14.135 3.220 ;
        RECT  13.715 2.520 13.975 3.220 ;
        END
        ANTENNAGATEAREA     0.3250 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.285 2.360 2.445 ;
        RECT  1.505 1.290 1.715 2.445 ;
        RECT  1.415 1.305 1.505 2.445 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.540 0.820 1.800 ;
        RECT  0.125 1.290 0.335 1.800 ;
        END
        ANTENNAGATEAREA     0.2652 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.900 1.700 6.320 2.095 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.295 0.595 16.455 2.320 ;
        RECT  14.795 0.595 16.295 0.755 ;
        RECT  15.510 2.160 16.295 2.320 ;
        RECT  15.510 2.520 15.515 3.220 ;
        RECT  15.305 2.160 15.510 3.220 ;
        RECT  15.240 2.160 15.305 3.100 ;
        RECT  14.535 0.595 14.795 1.195 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.115 1.290 17.355 2.745 ;
        RECT  16.895 1.290 17.115 1.450 ;
        RECT  16.520 2.505 17.115 2.745 ;
        RECT  16.795 1.105 16.895 1.450 ;
        RECT  16.635 0.645 16.795 1.450 ;
        RECT  16.260 2.505 16.520 3.105 ;
        RECT  16.225 2.745 16.260 2.995 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.700 2.175 1.990 ;
        RECT  1.895 1.530 2.150 2.085 ;
        END
        ANTENNAGATEAREA     0.2678 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.085 1.695 5.555 1.990 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.355 -0.250 17.480 0.250 ;
        RECT  17.095 -0.250 17.355 1.095 ;
        RECT  16.295 -0.250 17.095 0.250 ;
        RECT  16.035 -0.250 16.295 0.405 ;
        RECT  15.345 -0.250 16.035 0.250 ;
        RECT  15.085 -0.250 15.345 0.405 ;
        RECT  14.285 -0.250 15.085 0.250 ;
        RECT  14.025 -0.250 14.285 1.165 ;
        RECT  13.225 -0.250 14.025 0.250 ;
        RECT  12.965 -0.250 13.225 1.135 ;
        RECT  5.785 -0.250 12.965 0.250 ;
        RECT  5.525 -0.250 5.785 0.405 ;
        RECT  4.615 -0.250 5.525 0.250 ;
        RECT  4.355 -0.250 4.615 0.405 ;
        RECT  2.175 -0.250 4.355 0.250 ;
        RECT  1.915 -0.250 2.175 0.405 ;
        RECT  0.405 -0.250 1.915 0.250 ;
        RECT  0.145 -0.250 0.405 0.405 ;
        RECT  0.000 -0.250 0.145 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.045 3.440 17.480 3.940 ;
        RECT  16.785 2.955 17.045 3.940 ;
        RECT  16.010 3.440 16.785 3.940 ;
        RECT  15.750 2.600 16.010 3.940 ;
        RECT  14.965 3.440 15.750 3.940 ;
        RECT  14.705 2.445 14.965 3.940 ;
        RECT  11.750 3.440 14.705 3.940 ;
        RECT  11.150 3.285 11.750 3.940 ;
        RECT  8.440 3.440 11.150 3.940 ;
        RECT  8.180 3.105 8.440 3.940 ;
        RECT  6.930 3.440 8.180 3.940 ;
        RECT  5.990 3.050 6.930 3.940 ;
        RECT  4.470 3.440 5.990 3.940 ;
        RECT  4.210 3.285 4.470 3.940 ;
        RECT  2.105 3.440 4.210 3.940 ;
        RECT  1.845 3.005 2.105 3.940 ;
        RECT  0.385 3.440 1.845 3.940 ;
        RECT  0.125 2.555 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.940 0.955 16.100 1.980 ;
        RECT  15.485 0.955 15.940 1.115 ;
        RECT  15.055 1.820 15.940 1.980 ;
        RECT  14.525 1.470 15.645 1.630 ;
        RECT  14.895 1.820 15.055 2.265 ;
        RECT  14.415 2.105 14.895 2.265 ;
        RECT  14.365 1.470 14.525 1.920 ;
        RECT  14.155 2.105 14.415 2.740 ;
        RECT  12.400 1.760 14.365 1.920 ;
        RECT  13.340 2.105 14.155 2.265 ;
        RECT  13.515 0.555 13.775 1.580 ;
        RECT  13.275 2.780 13.535 3.105 ;
        RECT  12.765 1.420 13.515 1.580 ;
        RECT  13.080 2.105 13.340 2.365 ;
        RECT  8.990 2.945 13.275 3.105 ;
        RECT  12.645 2.505 12.805 2.765 ;
        RECT  12.605 0.480 12.765 1.580 ;
        RECT  9.395 2.605 12.645 2.765 ;
        RECT  12.490 0.480 12.605 0.640 ;
        RECT  12.230 0.470 12.490 0.640 ;
        RECT  12.400 2.245 12.450 2.405 ;
        RECT  12.240 0.875 12.400 2.405 ;
        RECT  10.675 0.875 12.240 1.035 ;
        RECT  10.110 2.245 12.240 2.405 ;
        RECT  8.860 0.480 12.230 0.640 ;
        RECT  11.720 1.215 11.980 1.545 ;
        RECT  10.360 1.215 11.720 1.375 ;
        RECT  11.265 1.555 11.525 1.765 ;
        RECT  9.930 1.605 11.265 1.765 ;
        RECT  10.200 0.820 10.360 1.375 ;
        RECT  9.305 0.820 10.200 0.980 ;
        RECT  9.770 1.160 9.930 2.245 ;
        RECT  9.665 1.160 9.770 1.320 ;
        RECT  8.635 2.085 9.770 2.245 ;
        RECT  9.305 1.560 9.590 1.830 ;
        RECT  9.235 2.425 9.395 2.765 ;
        RECT  9.145 0.820 9.305 1.830 ;
        RECT  7.245 2.425 9.235 2.585 ;
        RECT  8.515 0.940 9.145 1.100 ;
        RECT  8.830 2.765 8.990 3.105 ;
        RECT  8.700 0.480 8.860 0.755 ;
        RECT  8.730 2.765 8.830 2.940 ;
        RECT  7.890 2.765 8.730 2.925 ;
        RECT  8.475 1.335 8.635 2.245 ;
        RECT  8.355 0.585 8.515 1.100 ;
        RECT  8.175 1.335 8.475 1.495 ;
        RECT  7.080 2.085 8.475 2.245 ;
        RECT  5.195 0.585 8.355 0.745 ;
        RECT  7.970 1.675 8.235 1.890 ;
        RECT  8.015 0.925 8.175 1.495 ;
        RECT  7.915 0.925 8.015 1.185 ;
        RECT  6.660 1.730 7.970 1.890 ;
        RECT  7.165 1.025 7.915 1.185 ;
        RECT  7.620 2.765 7.890 2.940 ;
        RECT  7.085 2.425 7.245 2.870 ;
        RECT  6.900 0.925 7.165 1.185 ;
        RECT  5.655 2.710 7.085 2.870 ;
        RECT  4.485 0.925 6.900 1.085 ;
        RECT  6.660 2.365 6.770 2.525 ;
        RECT  6.500 1.280 6.660 2.525 ;
        RECT  6.125 1.280 6.500 1.440 ;
        RECT  5.495 2.170 5.655 2.910 ;
        RECT  4.825 2.170 5.495 2.330 ;
        RECT  5.300 3.100 5.440 3.260 ;
        RECT  5.140 2.510 5.300 3.260 ;
        RECT  4.825 1.275 5.215 1.435 ;
        RECT  4.935 0.540 5.195 0.745 ;
        RECT  3.805 2.510 5.140 2.670 ;
        RECT  4.800 2.850 4.960 3.110 ;
        RECT  3.415 0.585 4.935 0.745 ;
        RECT  4.665 1.275 4.825 2.330 ;
        RECT  3.925 2.850 4.800 3.010 ;
        RECT  4.635 1.695 4.665 2.330 ;
        RECT  4.145 1.695 4.635 1.855 ;
        RECT  4.325 0.925 4.485 1.425 ;
        RECT  4.225 1.165 4.325 1.425 ;
        RECT  3.985 1.650 4.145 1.910 ;
        RECT  3.715 2.850 3.925 3.045 ;
        RECT  3.645 0.925 3.805 2.670 ;
        RECT  3.330 2.885 3.715 3.045 ;
        RECT  3.595 0.925 3.645 1.185 ;
        RECT  3.510 2.270 3.645 2.670 ;
        RECT  3.415 1.330 3.465 1.590 ;
        RECT  3.330 0.585 3.415 1.590 ;
        RECT  3.255 0.585 3.330 3.045 ;
        RECT  3.170 1.330 3.255 3.045 ;
        RECT  2.990 0.495 3.075 1.095 ;
        RECT  2.915 0.495 2.990 3.060 ;
        RECT  2.830 0.585 2.915 3.060 ;
        RECT  1.315 0.585 2.830 0.745 ;
        RECT  1.275 2.645 2.830 2.805 ;
        RECT  2.460 0.950 2.620 2.000 ;
        RECT  1.170 0.950 2.460 1.110 ;
        RECT  1.055 0.510 1.315 0.770 ;
        RECT  1.015 2.605 1.275 3.205 ;
        RECT  1.010 0.950 1.170 2.155 ;
        RECT  0.635 0.950 1.010 1.295 ;
        RECT  0.875 1.995 1.010 2.155 ;
        RECT  0.615 1.995 0.875 2.255 ;
    END
END SDFFNSRX4

MACRO SDFFNSRX2
    CLASS CORE ;
    FOREIGN SDFFNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.230 2.785 10.575 3.220 ;
        END
        ANTENNAGATEAREA     0.1807 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.530 1.295 1.990 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.190 1.685 5.620 1.990 ;
        RECT  5.185 1.700 5.190 1.990 ;
        END
        ANTENNAGATEAREA     0.0650 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.280 2.110 12.295 2.400 ;
        RECT  12.120 0.620 12.280 2.400 ;
        RECT  12.085 0.620 12.120 0.945 ;
        RECT  12.085 2.110 12.120 2.400 ;
        RECT  11.190 0.620 12.085 0.780 ;
        RECT  11.845 2.240 12.085 2.400 ;
        RECT  11.585 2.240 11.845 2.510 ;
        RECT  11.145 0.565 11.190 0.780 ;
        RECT  10.885 0.565 11.145 1.165 ;
        END
        ANTENNADIFFAREA     0.6592 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.740 0.695 12.755 3.025 ;
        RECT  12.495 0.645 12.740 3.025 ;
        RECT  12.480 0.645 12.495 1.245 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.240 1.720 2.405 ;
        RECT  1.685 2.110 1.715 2.405 ;
        RECT  1.525 1.265 1.685 2.405 ;
        RECT  1.505 2.110 1.525 2.405 ;
        RECT  1.475 2.205 1.505 2.405 ;
        RECT  1.215 2.205 1.475 2.465 ;
        END
        ANTENNAGATEAREA     0.1430 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 1.695 4.935 1.990 ;
        END
        ANTENNAGATEAREA     0.0650 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.190 -0.250 12.880 0.250 ;
        RECT  11.930 -0.250 12.190 0.405 ;
        RECT  10.635 -0.250 11.930 0.250 ;
        RECT  10.375 -0.250 10.635 1.165 ;
        RECT  5.215 -0.250 10.375 0.250 ;
        RECT  4.955 -0.250 5.215 0.405 ;
        RECT  4.040 -0.250 4.955 0.250 ;
        RECT  3.780 -0.250 4.040 0.405 ;
        RECT  1.540 -0.250 3.780 0.250 ;
        RECT  1.280 -0.250 1.540 0.405 ;
        RECT  0.265 -0.250 1.280 0.250 ;
        RECT  0.265 1.035 0.385 1.295 ;
        RECT  0.105 -0.250 0.265 1.295 ;
        RECT  0.000 -0.250 0.105 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.245 3.440 12.880 3.940 ;
        RECT  11.985 2.935 12.245 3.940 ;
        RECT  11.335 3.440 11.985 3.940 ;
        RECT  11.075 2.185 11.335 3.940 ;
        RECT  8.565 3.440 11.075 3.940 ;
        RECT  8.305 3.105 8.565 3.940 ;
        RECT  7.045 3.440 8.305 3.940 ;
        RECT  6.785 3.105 7.045 3.940 ;
        RECT  5.845 3.440 6.785 3.940 ;
        RECT  5.585 3.105 5.845 3.940 ;
        RECT  4.035 3.440 5.585 3.940 ;
        RECT  3.775 3.285 4.035 3.940 ;
        RECT  1.675 3.440 3.775 3.940 ;
        RECT  1.415 3.285 1.675 3.940 ;
        RECT  0.385 3.440 1.415 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.885 1.605 11.935 1.865 ;
        RECT  11.725 0.965 11.885 2.005 ;
        RECT  11.395 0.965 11.725 1.125 ;
        RECT  10.670 1.845 11.725 2.005 ;
        RECT  10.885 1.350 11.485 1.645 ;
        RECT  10.090 1.350 10.885 1.510 ;
        RECT  10.570 1.845 10.670 2.485 ;
        RECT  10.410 1.745 10.570 2.485 ;
        RECT  9.670 1.745 10.410 1.905 ;
        RECT  9.865 0.475 10.125 1.075 ;
        RECT  9.930 1.275 10.090 1.510 ;
        RECT  9.890 2.085 10.050 3.085 ;
        RECT  9.390 1.275 9.930 1.435 ;
        RECT  9.190 2.085 9.890 2.245 ;
        RECT  8.920 2.925 9.890 3.085 ;
        RECT  9.790 0.475 9.865 0.635 ;
        RECT  9.630 0.455 9.790 0.635 ;
        RECT  9.550 2.425 9.710 2.745 ;
        RECT  9.410 1.645 9.670 1.905 ;
        RECT  9.005 0.455 9.630 0.615 ;
        RECT  7.595 2.425 9.550 2.585 ;
        RECT  9.185 0.795 9.445 0.975 ;
        RECT  9.230 1.165 9.390 1.435 ;
        RECT  8.680 1.165 9.230 1.325 ;
        RECT  9.030 1.735 9.190 2.245 ;
        RECT  8.340 0.815 9.185 0.975 ;
        RECT  9.020 1.735 9.030 1.895 ;
        RECT  8.860 1.635 9.020 1.895 ;
        RECT  8.845 0.455 9.005 0.630 ;
        RECT  8.760 2.765 8.920 3.085 ;
        RECT  7.120 0.470 8.845 0.630 ;
        RECT  8.680 2.085 8.845 2.245 ;
        RECT  5.245 2.765 8.760 2.925 ;
        RECT  8.520 1.165 8.680 2.245 ;
        RECT  8.180 0.815 8.340 1.785 ;
        RECT  7.955 1.965 8.215 2.245 ;
        RECT  7.480 0.815 8.180 0.975 ;
        RECT  8.080 1.525 8.180 1.785 ;
        RECT  7.900 1.165 7.965 1.325 ;
        RECT  7.900 1.965 7.955 2.125 ;
        RECT  7.740 1.165 7.900 2.125 ;
        RECT  7.705 1.165 7.740 1.445 ;
        RECT  6.440 1.285 7.705 1.445 ;
        RECT  7.335 2.305 7.595 2.585 ;
        RECT  7.320 0.815 7.480 1.100 ;
        RECT  6.590 2.425 7.335 2.585 ;
        RECT  6.780 0.940 7.320 1.100 ;
        RECT  6.960 0.470 7.120 0.755 ;
        RECT  6.620 0.545 6.780 1.100 ;
        RECT  6.040 0.545 6.620 0.705 ;
        RECT  6.430 1.865 6.590 2.585 ;
        RECT  6.280 0.885 6.440 1.445 ;
        RECT  6.310 1.865 6.430 2.125 ;
        RECT  3.920 0.925 6.280 1.085 ;
        RECT  5.985 2.425 6.245 2.585 ;
        RECT  5.985 1.405 6.100 1.665 ;
        RECT  5.880 0.545 6.040 0.745 ;
        RECT  5.825 1.265 5.985 2.585 ;
        RECT  2.850 0.585 5.880 0.745 ;
        RECT  5.390 1.265 5.825 1.425 ;
        RECT  5.085 2.170 5.245 2.925 ;
        RECT  4.285 2.170 5.085 2.330 ;
        RECT  4.905 3.100 5.005 3.260 ;
        RECT  4.745 2.510 4.905 3.260 ;
        RECT  3.190 2.510 4.745 2.670 ;
        RECT  4.285 1.265 4.615 1.425 ;
        RECT  4.405 2.850 4.565 3.110 ;
        RECT  3.440 2.850 4.405 3.010 ;
        RECT  4.125 1.265 4.285 2.330 ;
        RECT  3.530 1.645 4.125 1.805 ;
        RECT  3.760 0.925 3.920 1.435 ;
        RECT  3.660 1.175 3.760 1.435 ;
        RECT  3.370 1.645 3.530 1.915 ;
        RECT  3.180 2.850 3.440 3.110 ;
        RECT  3.030 0.925 3.190 2.670 ;
        RECT  2.850 2.850 3.180 3.010 ;
        RECT  2.815 0.585 2.850 3.010 ;
        RECT  2.690 0.535 2.815 3.010 ;
        RECT  2.555 0.535 2.690 0.745 ;
        RECT  2.370 0.965 2.510 2.875 ;
        RECT  2.350 0.585 2.370 2.875 ;
        RECT  2.210 0.585 2.350 1.125 ;
        RECT  2.225 2.275 2.350 2.875 ;
        RECT  0.825 2.645 2.225 2.805 ;
        RECT  0.605 0.585 2.210 0.745 ;
        RECT  2.030 1.410 2.170 1.670 ;
        RECT  1.870 0.925 2.030 1.670 ;
        RECT  0.970 0.925 1.870 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.665 0.925 0.825 2.215 ;
        RECT  0.565 2.645 0.825 2.905 ;
        RECT  0.445 0.455 0.605 0.745 ;
    END
END SDFFNSRX2

MACRO SDFFNSRX1
    CLASS CORE ;
    FOREIGN SDFFNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 2.520 10.455 2.810 ;
        RECT  10.245 2.520 10.405 3.005 ;
        RECT  9.890 2.845 10.245 3.005 ;
        RECT  9.630 2.845 9.890 3.105 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.480 1.255 2.045 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.1105 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 1.700 5.725 1.960 ;
        RECT  5.370 1.290 5.395 1.960 ;
        RECT  5.235 1.290 5.370 1.860 ;
        RECT  5.185 1.290 5.235 1.765 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.230 0.645 11.390 2.925 ;
        RECT  11.165 0.645 11.230 0.945 ;
        RECT  11.165 2.335 11.230 2.925 ;
        RECT  10.920 0.645 11.165 0.805 ;
        RECT  10.920 2.765 11.165 2.925 ;
        RECT  10.660 0.545 10.920 0.805 ;
        RECT  10.660 2.765 10.920 3.025 ;
        END
        ANTENNADIFFAREA     0.3922 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.830 1.105 11.835 2.590 ;
        RECT  11.625 0.920 11.830 2.750 ;
        RECT  11.570 0.920 11.625 1.180 ;
        RECT  11.570 2.150 11.625 2.750 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.695 1.270 1.715 2.400 ;
        RECT  1.505 1.270 1.695 2.535 ;
        RECT  1.445 1.270 1.505 1.530 ;
        RECT  1.215 2.275 1.505 2.535 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.610 1.625 5.005 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.430 -0.250 11.960 0.250 ;
        RECT  11.170 -0.250 11.430 0.405 ;
        RECT  10.350 -0.250 11.170 0.250 ;
        RECT  10.090 -0.250 10.350 1.135 ;
        RECT  6.495 -0.250 10.090 0.250 ;
        RECT  5.895 -0.250 6.495 0.405 ;
        RECT  3.980 -0.250 5.895 0.250 ;
        RECT  3.720 -0.250 3.980 0.405 ;
        RECT  1.675 -0.250 3.720 0.250 ;
        RECT  1.415 -0.250 1.675 0.405 ;
        RECT  0.275 -0.250 1.415 0.250 ;
        RECT  0.275 1.035 0.335 1.295 ;
        RECT  0.115 -0.250 0.275 1.295 ;
        RECT  0.000 -0.250 0.115 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.430 3.440 11.960 3.940 ;
        RECT  11.170 3.285 11.430 3.940 ;
        RECT  10.350 3.440 11.170 3.940 ;
        RECT  10.090 3.285 10.350 3.940 ;
        RECT  8.265 3.440 10.090 3.940 ;
        RECT  8.005 3.115 8.265 3.940 ;
        RECT  6.545 3.440 8.005 3.940 ;
        RECT  5.605 3.055 6.545 3.940 ;
        RECT  4.045 3.440 5.605 3.940 ;
        RECT  3.785 3.285 4.045 3.940 ;
        RECT  1.675 3.440 3.785 3.940 ;
        RECT  1.415 3.285 1.675 3.940 ;
        RECT  0.385 3.440 1.415 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.945 1.635 11.050 1.895 ;
        RECT  10.785 1.120 10.945 2.345 ;
        RECT  10.660 1.120 10.785 1.380 ;
        RECT  10.660 2.065 10.785 2.345 ;
        RECT  9.555 2.065 10.660 2.225 ;
        RECT  10.200 1.510 10.460 1.770 ;
        RECT  9.345 1.530 10.200 1.690 ;
        RECT  9.710 0.805 9.810 1.065 ;
        RECT  9.495 2.405 9.755 2.665 ;
        RECT  9.550 0.470 9.710 1.065 ;
        RECT  9.295 1.965 9.555 2.225 ;
        RECT  7.085 0.470 9.550 0.630 ;
        RECT  9.380 2.505 9.495 2.665 ;
        RECT  9.220 2.505 9.380 2.935 ;
        RECT  9.185 1.250 9.345 1.690 ;
        RECT  7.090 2.775 9.220 2.935 ;
        RECT  8.665 1.250 9.185 1.410 ;
        RECT  8.870 0.810 9.130 1.070 ;
        RECT  8.845 1.655 9.005 2.595 ;
        RECT  8.225 0.810 8.870 0.970 ;
        RECT  8.745 1.655 8.845 1.915 ;
        RECT  7.430 2.435 8.845 2.595 ;
        RECT  8.565 1.150 8.665 1.410 ;
        RECT  8.565 2.095 8.665 2.255 ;
        RECT  8.405 1.150 8.565 2.255 ;
        RECT  8.065 0.810 8.225 2.050 ;
        RECT  7.425 0.810 8.065 0.970 ;
        RECT  7.785 2.095 7.885 2.255 ;
        RECT  7.785 1.150 7.865 1.310 ;
        RECT  7.625 1.150 7.785 2.255 ;
        RECT  7.605 1.150 7.625 1.625 ;
        RECT  6.405 1.465 7.605 1.625 ;
        RECT  7.270 2.160 7.430 2.595 ;
        RECT  7.265 0.810 7.425 1.285 ;
        RECT  6.650 2.160 7.270 2.320 ;
        RECT  6.745 1.125 7.265 1.285 ;
        RECT  6.830 2.515 7.090 2.935 ;
        RECT  6.925 0.470 7.085 0.945 ;
        RECT  6.065 1.805 6.920 1.965 ;
        RECT  6.585 0.585 6.745 1.285 ;
        RECT  6.490 2.160 6.650 2.805 ;
        RECT  5.685 0.585 6.585 0.745 ;
        RECT  5.245 2.645 6.490 2.805 ;
        RECT  6.245 0.925 6.405 1.625 ;
        RECT  5.345 0.925 6.245 1.085 ;
        RECT  5.905 1.265 6.065 2.465 ;
        RECT  5.805 1.265 5.905 1.425 ;
        RECT  5.705 2.205 5.905 2.465 ;
        RECT  5.525 0.470 5.685 0.745 ;
        RECT  4.625 0.470 5.525 0.630 ;
        RECT  5.185 0.845 5.345 1.085 ;
        RECT  5.085 2.170 5.245 2.910 ;
        RECT  4.665 0.845 5.185 1.005 ;
        RECT  4.430 2.170 5.085 2.330 ;
        RECT  4.905 3.100 5.085 3.260 ;
        RECT  4.845 1.185 5.005 1.445 ;
        RECT  4.745 2.510 4.905 3.260 ;
        RECT  4.430 1.285 4.845 1.445 ;
        RECT  3.185 2.510 4.745 2.670 ;
        RECT  4.505 0.845 4.665 1.085 ;
        RECT  4.365 0.445 4.625 0.630 ;
        RECT  4.405 2.850 4.565 3.110 ;
        RECT  3.985 0.925 4.505 1.085 ;
        RECT  4.270 1.285 4.430 2.330 ;
        RECT  3.435 2.850 4.405 3.010 ;
        RECT  4.325 0.470 4.365 0.630 ;
        RECT  4.165 0.470 4.325 0.745 ;
        RECT  3.625 1.645 4.270 1.805 ;
        RECT  4.225 2.170 4.270 2.330 ;
        RECT  2.845 0.585 4.165 0.745 ;
        RECT  3.825 0.925 3.985 1.425 ;
        RECT  3.725 1.165 3.825 1.425 ;
        RECT  3.365 1.645 3.625 1.910 ;
        RECT  3.175 2.850 3.435 3.110 ;
        RECT  3.185 0.925 3.205 1.185 ;
        RECT  3.025 0.925 3.185 2.670 ;
        RECT  2.845 2.850 3.175 3.010 ;
        RECT  2.685 0.585 2.845 3.010 ;
        RECT  2.345 0.520 2.505 2.905 ;
        RECT  0.715 0.585 2.345 0.745 ;
        RECT  0.745 2.745 2.345 2.905 ;
        RECT  1.975 0.925 2.135 1.715 ;
        RECT  0.970 0.925 1.975 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.665 0.925 0.825 2.305 ;
        RECT  0.485 2.645 0.745 2.905 ;
        RECT  0.455 0.440 0.715 0.745 ;
    END
END SDFFNSRX1

MACRO SDFFNSRXL
    CLASS CORE ;
    FOREIGN SDFFNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 2.520 10.455 2.810 ;
        RECT  10.245 2.520 10.405 3.005 ;
        RECT  9.890 2.845 10.245 3.005 ;
        RECT  9.630 2.845 9.890 3.105 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.475 1.295 2.065 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.565 1.700 5.725 2.025 ;
        RECT  5.395 1.700 5.565 1.990 ;
        RECT  5.370 1.290 5.395 1.990 ;
        RECT  5.235 1.290 5.370 1.860 ;
        RECT  5.185 1.290 5.235 1.765 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.230 0.645 11.390 2.925 ;
        RECT  11.165 0.645 11.230 0.945 ;
        RECT  11.165 2.335 11.230 2.925 ;
        RECT  10.890 0.645 11.165 0.805 ;
        RECT  10.920 2.765 11.165 2.925 ;
        RECT  10.660 2.765 10.920 3.025 ;
        RECT  10.630 0.545 10.890 0.805 ;
        END
        ANTENNADIFFAREA     0.2231 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.830 1.105 11.835 2.185 ;
        RECT  11.625 0.920 11.830 2.580 ;
        RECT  11.570 0.920 11.625 1.180 ;
        RECT  11.570 2.320 11.625 2.580 ;
        END
        ANTENNADIFFAREA     0.2135 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.265 1.735 1.525 ;
        RECT  1.505 1.265 1.715 2.505 ;
        RECT  1.475 1.265 1.505 1.765 ;
        RECT  1.235 2.245 1.505 2.505 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 1.645 5.005 1.925 ;
        RECT  4.845 1.645 4.935 1.990 ;
        RECT  4.465 1.695 4.845 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.400 -0.250 11.960 0.250 ;
        RECT  11.140 -0.250 11.400 0.405 ;
        RECT  10.320 -0.250 11.140 0.250 ;
        RECT  10.060 -0.250 10.320 1.135 ;
        RECT  6.495 -0.250 10.060 0.250 ;
        RECT  5.895 -0.250 6.495 0.405 ;
        RECT  3.980 -0.250 5.895 0.250 ;
        RECT  3.720 -0.250 3.980 0.405 ;
        RECT  1.605 -0.250 3.720 0.250 ;
        RECT  1.345 -0.250 1.605 0.405 ;
        RECT  0.285 -0.250 1.345 0.250 ;
        RECT  0.285 1.035 0.385 1.295 ;
        RECT  0.125 -0.250 0.285 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.430 3.440 11.960 3.940 ;
        RECT  11.170 3.285 11.430 3.940 ;
        RECT  10.350 3.440 11.170 3.940 ;
        RECT  10.090 3.285 10.350 3.940 ;
        RECT  8.265 3.440 10.090 3.940 ;
        RECT  8.005 3.115 8.265 3.940 ;
        RECT  6.545 3.440 8.005 3.940 ;
        RECT  5.605 3.055 6.545 3.940 ;
        RECT  4.045 3.440 5.605 3.940 ;
        RECT  3.785 3.285 4.045 3.940 ;
        RECT  1.675 3.440 3.785 3.940 ;
        RECT  1.415 3.285 1.675 3.940 ;
        RECT  0.385 3.440 1.415 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.950 1.635 11.050 1.895 ;
        RECT  10.790 1.120 10.950 2.345 ;
        RECT  10.630 1.120 10.790 1.380 ;
        RECT  10.660 2.085 10.790 2.345 ;
        RECT  10.215 2.135 10.660 2.295 ;
        RECT  10.190 1.510 10.450 1.770 ;
        RECT  10.055 2.010 10.215 2.295 ;
        RECT  9.735 1.510 10.190 1.670 ;
        RECT  9.550 2.010 10.055 2.170 ;
        RECT  9.680 0.695 9.780 0.955 ;
        RECT  9.490 2.405 9.750 2.665 ;
        RECT  9.575 1.315 9.735 1.670 ;
        RECT  9.520 0.470 9.680 0.955 ;
        RECT  8.660 1.315 9.575 1.475 ;
        RECT  9.290 1.910 9.550 2.170 ;
        RECT  7.085 0.470 9.520 0.630 ;
        RECT  9.380 2.505 9.490 2.665 ;
        RECT  9.220 2.505 9.380 2.935 ;
        RECT  7.090 2.775 9.220 2.935 ;
        RECT  8.840 0.810 9.100 1.135 ;
        RECT  8.850 1.655 9.010 2.595 ;
        RECT  8.745 1.655 8.850 1.915 ;
        RECT  7.435 2.435 8.850 2.595 ;
        RECT  8.220 0.810 8.840 0.970 ;
        RECT  8.560 2.095 8.665 2.255 ;
        RECT  8.560 1.150 8.660 1.475 ;
        RECT  8.400 1.150 8.560 2.255 ;
        RECT  8.060 0.810 8.220 2.050 ;
        RECT  7.425 0.810 8.060 0.970 ;
        RECT  7.775 2.095 7.875 2.255 ;
        RECT  7.775 1.150 7.865 1.310 ;
        RECT  7.615 1.150 7.775 2.255 ;
        RECT  7.605 1.150 7.615 1.610 ;
        RECT  6.405 1.450 7.605 1.610 ;
        RECT  7.275 2.230 7.435 2.595 ;
        RECT  7.265 0.810 7.425 1.270 ;
        RECT  6.545 2.230 7.275 2.390 ;
        RECT  6.745 1.110 7.265 1.270 ;
        RECT  6.830 2.570 7.090 2.935 ;
        RECT  6.925 0.470 7.085 0.925 ;
        RECT  6.660 1.790 6.920 2.050 ;
        RECT  6.585 0.585 6.745 1.270 ;
        RECT  6.065 1.890 6.660 2.050 ;
        RECT  5.685 0.585 6.585 0.745 ;
        RECT  6.385 2.230 6.545 2.830 ;
        RECT  6.245 0.925 6.405 1.610 ;
        RECT  5.245 2.670 6.385 2.830 ;
        RECT  5.345 0.925 6.245 1.085 ;
        RECT  5.905 1.265 6.065 2.465 ;
        RECT  5.805 1.265 5.905 1.425 ;
        RECT  5.705 2.205 5.905 2.465 ;
        RECT  5.525 0.470 5.685 0.745 ;
        RECT  4.625 0.470 5.525 0.630 ;
        RECT  5.185 0.845 5.345 1.085 ;
        RECT  5.085 2.170 5.245 2.910 ;
        RECT  4.665 0.845 5.185 1.005 ;
        RECT  4.905 3.100 5.185 3.260 ;
        RECT  4.285 2.170 5.085 2.330 ;
        RECT  4.845 1.185 5.005 1.445 ;
        RECT  4.745 2.510 4.905 3.260 ;
        RECT  4.285 1.285 4.845 1.445 ;
        RECT  3.185 2.510 4.745 2.670 ;
        RECT  4.505 0.845 4.665 1.085 ;
        RECT  4.365 0.445 4.625 0.630 ;
        RECT  4.405 2.850 4.565 3.110 ;
        RECT  3.935 0.925 4.505 1.085 ;
        RECT  3.435 2.850 4.405 3.010 ;
        RECT  4.325 0.470 4.365 0.630 ;
        RECT  4.165 0.470 4.325 0.745 ;
        RECT  4.125 1.285 4.285 2.330 ;
        RECT  2.845 0.585 4.165 0.745 ;
        RECT  3.625 1.650 4.125 1.810 ;
        RECT  3.775 0.925 3.935 1.425 ;
        RECT  3.675 1.165 3.775 1.425 ;
        RECT  3.365 1.650 3.625 1.910 ;
        RECT  3.175 2.850 3.435 3.110 ;
        RECT  3.025 0.925 3.185 2.670 ;
        RECT  2.845 2.850 3.175 3.010 ;
        RECT  2.685 0.585 2.845 3.010 ;
        RECT  2.345 0.455 2.505 2.905 ;
        RECT  0.725 0.585 2.345 0.745 ;
        RECT  0.745 2.745 2.345 2.905 ;
        RECT  2.005 0.925 2.165 1.715 ;
        RECT  0.970 0.925 2.005 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.665 0.925 0.825 2.305 ;
        RECT  0.485 2.645 0.745 2.905 ;
        RECT  0.465 0.440 0.725 0.745 ;
    END
END SDFFNSRXL

MACRO SDFFSRX4
    CLASS CORE ;
    FOREIGN SDFFSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.960 2.930 14.135 3.220 ;
        RECT  13.800 2.505 13.960 3.220 ;
        RECT  13.670 2.505 13.800 2.765 ;
        END
        ANTENNAGATEAREA     0.3250 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 2.260 2.295 2.420 ;
        RECT  1.255 1.320 1.505 1.480 ;
        RECT  1.095 1.320 1.255 2.420 ;
        RECT  1.045 1.515 1.095 2.175 ;
        END
        ANTENNAGATEAREA     0.1326 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.490 0.505 1.750 ;
        RECT  0.125 1.290 0.335 1.750 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.220 2.110 6.315 2.400 ;
        RECT  6.060 1.620 6.220 2.400 ;
        RECT  5.960 1.620 6.060 1.880 ;
        END
        ANTENNAGATEAREA     0.1144 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.290 0.595 16.450 2.345 ;
        RECT  14.795 0.595 16.290 0.755 ;
        RECT  15.515 2.185 16.290 2.345 ;
        RECT  15.305 2.185 15.515 3.220 ;
        RECT  15.240 2.185 15.305 3.125 ;
        RECT  14.535 0.595 14.795 1.195 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.160 1.290 17.355 1.990 ;
        RECT  17.145 1.085 17.160 1.990 ;
        RECT  16.795 1.085 17.145 2.765 ;
        RECT  16.685 0.645 16.795 2.765 ;
        RECT  16.635 0.645 16.685 1.245 ;
        RECT  16.520 2.525 16.685 2.765 ;
        RECT  16.260 2.525 16.520 3.125 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.760 1.600 2.020 1.860 ;
        RECT  1.715 1.700 1.760 1.860 ;
        RECT  1.505 1.700 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.2717 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 1.645 5.395 1.860 ;
        RECT  4.475 1.700 5.135 1.860 ;
        RECT  4.265 1.700 4.475 1.990 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.355 -0.250 17.480 0.250 ;
        RECT  17.095 -0.250 17.355 0.795 ;
        RECT  16.295 -0.250 17.095 0.250 ;
        RECT  16.035 -0.250 16.295 0.405 ;
        RECT  15.345 -0.250 16.035 0.250 ;
        RECT  15.085 -0.250 15.345 0.405 ;
        RECT  14.285 -0.250 15.085 0.250 ;
        RECT  14.025 -0.250 14.285 1.165 ;
        RECT  13.225 -0.250 14.025 0.250 ;
        RECT  12.965 -0.250 13.225 1.135 ;
        RECT  5.785 -0.250 12.965 0.250 ;
        RECT  5.525 -0.250 5.785 0.405 ;
        RECT  4.505 -0.250 5.525 0.250 ;
        RECT  4.245 -0.250 4.505 0.405 ;
        RECT  2.065 -0.250 4.245 0.250 ;
        RECT  1.805 -0.250 2.065 0.405 ;
        RECT  0.385 -0.250 1.805 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.045 3.440 17.480 3.940 ;
        RECT  16.785 2.955 17.045 3.940 ;
        RECT  16.010 3.440 16.785 3.940 ;
        RECT  15.750 2.600 16.010 3.940 ;
        RECT  14.965 3.440 15.750 3.940 ;
        RECT  14.705 2.445 14.965 3.940 ;
        RECT  11.720 3.440 14.705 3.940 ;
        RECT  11.120 3.285 11.720 3.940 ;
        RECT  8.440 3.440 11.120 3.940 ;
        RECT  8.180 3.105 8.440 3.940 ;
        RECT  6.920 3.440 8.180 3.940 ;
        RECT  5.980 3.105 6.920 3.940 ;
        RECT  4.410 3.440 5.980 3.940 ;
        RECT  4.150 3.080 4.410 3.940 ;
        RECT  2.035 3.440 4.150 3.940 ;
        RECT  1.775 2.955 2.035 3.940 ;
        RECT  0.385 3.440 1.775 3.940 ;
        RECT  0.125 2.480 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.940 0.955 16.100 2.005 ;
        RECT  15.485 0.955 15.940 1.115 ;
        RECT  15.890 1.605 15.940 2.005 ;
        RECT  14.415 1.845 15.890 2.005 ;
        RECT  14.365 1.405 15.645 1.665 ;
        RECT  14.255 1.845 14.415 2.710 ;
        RECT  14.075 1.505 14.365 1.665 ;
        RECT  14.155 2.145 14.255 2.710 ;
        RECT  13.320 2.145 14.155 2.305 ;
        RECT  13.915 1.505 14.075 1.815 ;
        RECT  12.415 1.655 13.915 1.815 ;
        RECT  13.675 0.645 13.775 1.245 ;
        RECT  13.515 0.645 13.675 1.475 ;
        RECT  13.260 2.945 13.520 3.230 ;
        RECT  12.765 1.315 13.515 1.475 ;
        RECT  13.060 2.080 13.320 2.340 ;
        RECT  8.990 2.945 13.260 3.105 ;
        RECT  12.630 2.500 12.790 2.765 ;
        RECT  12.605 0.470 12.765 1.475 ;
        RECT  9.415 2.605 12.630 2.765 ;
        RECT  9.930 0.470 12.605 0.630 ;
        RECT  12.415 2.265 12.450 2.425 ;
        RECT  12.255 0.815 12.415 2.425 ;
        RECT  10.670 0.815 12.255 0.975 ;
        RECT  10.245 2.265 12.255 2.425 ;
        RECT  11.910 1.160 12.070 2.085 ;
        RECT  9.735 1.160 11.910 1.320 ;
        RECT  10.720 1.925 11.910 2.085 ;
        RECT  11.470 1.535 11.730 1.725 ;
        RECT  8.870 1.535 11.470 1.695 ;
        RECT  10.560 1.890 10.720 2.085 ;
        RECT  9.540 1.890 10.560 2.050 ;
        RECT  9.985 2.245 10.245 2.425 ;
        RECT  9.670 0.470 9.930 0.735 ;
        RECT  9.575 0.925 9.735 1.320 ;
        RECT  8.910 0.470 9.670 0.630 ;
        RECT  8.350 0.925 9.575 1.085 ;
        RECT  9.380 1.890 9.540 2.245 ;
        RECT  9.255 2.425 9.415 2.765 ;
        RECT  7.080 2.085 9.380 2.245 ;
        RECT  7.265 2.425 9.255 2.585 ;
        RECT  8.730 2.765 8.990 3.105 ;
        RECT  8.650 0.470 8.910 0.745 ;
        RECT  8.710 1.265 8.870 1.695 ;
        RECT  7.890 2.765 8.730 2.925 ;
        RECT  6.900 1.265 8.710 1.425 ;
        RECT  8.090 0.825 8.350 1.085 ;
        RECT  7.970 1.645 8.230 1.905 ;
        RECT  7.340 0.925 8.090 1.085 ;
        RECT  6.710 1.745 7.970 1.905 ;
        RECT  7.620 2.765 7.890 2.940 ;
        RECT  7.240 0.825 7.340 1.085 ;
        RECT  7.105 2.425 7.265 2.875 ;
        RECT  7.080 0.595 7.240 1.085 ;
        RECT  5.100 2.715 7.105 2.875 ;
        RECT  5.430 0.595 7.080 0.755 ;
        RECT  6.740 0.935 6.900 1.425 ;
        RECT  6.710 2.355 6.820 2.515 ;
        RECT  5.780 0.935 6.740 1.095 ;
        RECT  6.560 1.745 6.710 2.515 ;
        RECT  6.550 1.275 6.560 2.515 ;
        RECT  6.400 1.275 6.550 1.910 ;
        RECT  6.125 1.275 6.400 1.435 ;
        RECT  5.620 0.935 5.780 2.535 ;
        RECT  4.955 1.275 5.620 1.435 ;
        RECT  5.440 2.325 5.620 2.535 ;
        RECT  4.755 3.060 5.550 3.220 ;
        RECT  5.280 2.045 5.440 2.535 ;
        RECT  5.270 0.595 5.430 1.090 ;
        RECT  4.655 2.045 5.280 2.205 ;
        RECT  4.405 0.930 5.270 1.090 ;
        RECT  4.940 2.390 5.100 2.875 ;
        RECT  3.820 0.585 5.085 0.745 ;
        RECT  4.070 2.390 4.940 2.550 ;
        RECT  4.595 2.735 4.755 3.220 ;
        RECT  3.510 2.735 4.595 2.895 ;
        RECT  4.245 0.930 4.405 1.515 ;
        RECT  4.145 1.255 4.245 1.515 ;
        RECT  3.910 1.750 4.070 2.550 ;
        RECT  3.820 1.750 3.910 1.910 ;
        RECT  3.660 0.470 3.820 1.910 ;
        RECT  3.490 0.470 3.660 0.630 ;
        RECT  3.390 1.650 3.660 1.910 ;
        RECT  3.250 2.120 3.510 3.105 ;
        RECT  3.380 0.865 3.480 1.125 ;
        RECT  3.220 0.865 3.380 1.465 ;
        RECT  3.190 2.120 3.250 2.280 ;
        RECT  3.190 1.305 3.220 1.465 ;
        RECT  3.030 1.305 3.190 2.280 ;
        RECT  2.850 2.470 2.975 3.070 ;
        RECT  2.850 0.510 2.970 1.110 ;
        RECT  2.715 0.510 2.850 3.070 ;
        RECT  2.710 0.510 2.715 2.765 ;
        RECT  2.690 0.585 2.710 2.765 ;
        RECT  1.185 0.585 2.690 0.745 ;
        RECT  1.215 2.605 2.690 2.765 ;
        RECT  2.400 1.730 2.500 1.990 ;
        RECT  2.240 0.925 2.400 1.990 ;
        RECT  0.855 0.925 2.240 1.085 ;
        RECT  0.955 2.605 1.215 3.215 ;
        RECT  0.925 0.485 1.185 0.745 ;
        RECT  0.695 0.925 0.855 2.215 ;
        RECT  0.555 0.925 0.695 1.295 ;
        RECT  0.555 1.955 0.695 2.215 ;
    END
END SDFFSRX4

MACRO SDFFSRX2
    CLASS CORE ;
    FOREIGN SDFFSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.250 2.785 10.525 3.220 ;
        RECT  10.245 2.930 10.250 3.220 ;
        RECT  10.230 2.960 10.245 3.220 ;
        END
        ANTENNAGATEAREA     0.1807 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.520 1.295 1.985 ;
        RECT  1.045 1.520 1.255 1.990 ;
        RECT  1.005 1.520 1.045 1.985 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.585 2.000 5.855 2.470 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.280 2.110 12.295 2.400 ;
        RECT  12.245 0.620 12.280 2.400 ;
        RECT  12.120 0.620 12.245 2.410 ;
        RECT  12.085 0.620 12.120 0.975 ;
        RECT  12.085 2.110 12.120 2.410 ;
        RECT  11.220 0.620 12.085 0.780 ;
        RECT  11.845 2.250 12.085 2.410 ;
        RECT  11.585 2.250 11.845 2.510 ;
        RECT  11.145 0.490 11.220 0.780 ;
        RECT  10.885 0.490 11.145 1.090 ;
        END
        ANTENNADIFFAREA     0.6592 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.495 0.595 12.755 3.025 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.690 2.110 1.715 2.465 ;
        RECT  1.530 1.395 1.690 2.465 ;
        RECT  1.505 2.110 1.530 2.465 ;
        RECT  1.215 2.205 1.505 2.465 ;
        END
        ANTENNAGATEAREA     0.1430 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 1.700 5.395 1.990 ;
        RECT  4.705 1.830 5.185 1.990 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.215 -0.250 12.880 0.250 ;
        RECT  11.955 -0.250 12.215 0.405 ;
        RECT  10.635 -0.250 11.955 0.250 ;
        RECT  10.375 -0.250 10.635 1.090 ;
        RECT  5.285 -0.250 10.375 0.250 ;
        RECT  5.025 -0.250 5.285 0.405 ;
        RECT  3.785 -0.250 5.025 0.250 ;
        RECT  3.525 -0.250 3.785 0.585 ;
        RECT  1.565 -0.250 3.525 0.250 ;
        RECT  1.305 -0.250 1.565 0.405 ;
        RECT  0.265 -0.250 1.305 0.250 ;
        RECT  0.265 1.035 0.385 1.295 ;
        RECT  0.105 -0.250 0.265 1.295 ;
        RECT  0.000 -0.250 0.105 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.245 3.440 12.880 3.940 ;
        RECT  11.985 2.935 12.245 3.940 ;
        RECT  11.335 3.440 11.985 3.940 ;
        RECT  11.075 2.185 11.335 3.940 ;
        RECT  8.565 3.440 11.075 3.940 ;
        RECT  8.305 3.115 8.565 3.940 ;
        RECT  7.045 3.440 8.305 3.940 ;
        RECT  6.785 3.115 7.045 3.940 ;
        RECT  5.500 3.440 6.785 3.940 ;
        RECT  4.895 3.115 5.500 3.940 ;
        RECT  1.675 3.440 4.895 3.940 ;
        RECT  1.415 3.285 1.675 3.940 ;
        RECT  0.385 3.440 1.415 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.905 1.605 11.935 1.940 ;
        RECT  11.745 0.965 11.905 1.940 ;
        RECT  11.395 0.965 11.745 1.125 ;
        RECT  10.755 1.780 11.745 1.940 ;
        RECT  11.215 1.305 11.485 1.595 ;
        RECT  10.885 1.270 11.215 1.595 ;
        RECT  10.090 1.270 10.885 1.430 ;
        RECT  10.655 1.780 10.755 2.485 ;
        RECT  10.495 1.620 10.655 2.485 ;
        RECT  9.410 1.620 10.495 1.780 ;
        RECT  9.865 0.490 10.125 1.090 ;
        RECT  9.930 1.270 10.090 1.440 ;
        RECT  9.890 1.960 10.050 3.025 ;
        RECT  9.215 1.280 9.930 1.440 ;
        RECT  9.190 1.960 9.890 2.120 ;
        RECT  9.340 2.865 9.890 3.025 ;
        RECT  9.790 0.490 9.865 0.650 ;
        RECT  9.630 0.465 9.790 0.650 ;
        RECT  9.550 2.300 9.710 2.595 ;
        RECT  9.000 0.465 9.630 0.625 ;
        RECT  7.595 2.435 9.550 2.595 ;
        RECT  9.185 0.805 9.445 0.975 ;
        RECT  9.180 2.775 9.340 3.025 ;
        RECT  8.955 1.175 9.215 1.440 ;
        RECT  9.030 1.735 9.190 2.120 ;
        RECT  8.305 0.815 9.185 0.975 ;
        RECT  6.605 2.775 9.180 2.935 ;
        RECT  9.020 1.735 9.030 1.895 ;
        RECT  8.860 1.635 9.020 1.895 ;
        RECT  8.840 0.465 9.000 0.630 ;
        RECT  8.665 1.280 8.955 1.440 ;
        RECT  8.665 2.095 8.845 2.255 ;
        RECT  7.120 0.470 8.840 0.630 ;
        RECT  8.505 1.280 8.665 2.255 ;
        RECT  8.145 0.815 8.305 1.890 ;
        RECT  7.965 2.095 8.215 2.255 ;
        RECT  7.520 0.815 8.145 0.975 ;
        RECT  7.805 1.165 7.965 2.255 ;
        RECT  7.705 1.165 7.805 1.480 ;
        RECT  6.440 1.315 7.705 1.480 ;
        RECT  7.335 2.305 7.595 2.595 ;
        RECT  7.360 0.815 7.520 1.135 ;
        RECT  6.780 0.975 7.360 1.135 ;
        RECT  6.635 2.435 7.335 2.595 ;
        RECT  6.960 0.470 7.120 0.795 ;
        RECT  6.620 0.540 6.780 1.135 ;
        RECT  6.475 1.865 6.635 2.595 ;
        RECT  6.085 0.540 6.620 0.700 ;
        RECT  6.445 2.775 6.605 2.980 ;
        RECT  6.425 1.865 6.475 2.125 ;
        RECT  5.855 2.820 6.445 2.980 ;
        RECT  6.280 0.885 6.440 1.480 ;
        RECT  5.005 0.925 6.280 1.085 ;
        RECT  6.100 1.660 6.225 2.640 ;
        RECT  6.065 1.265 6.100 2.640 ;
        RECT  5.925 0.540 6.085 0.745 ;
        RECT  5.940 1.265 6.065 1.820 ;
        RECT  6.035 2.375 6.065 2.640 ;
        RECT  5.840 1.265 5.940 1.555 ;
        RECT  4.655 0.585 5.925 0.745 ;
        RECT  5.695 2.775 5.855 2.980 ;
        RECT  5.455 1.265 5.840 1.505 ;
        RECT  4.615 2.775 5.695 2.935 ;
        RECT  4.885 2.235 5.145 2.585 ;
        RECT  4.845 0.925 5.005 1.640 ;
        RECT  4.485 2.235 4.885 2.395 ;
        RECT  4.005 1.480 4.845 1.640 ;
        RECT  4.495 0.585 4.655 1.300 ;
        RECT  4.355 2.575 4.615 2.935 ;
        RECT  3.560 1.110 4.495 1.270 ;
        RECT  4.225 2.135 4.485 2.395 ;
        RECT  3.540 2.575 4.355 2.735 ;
        RECT  4.155 0.530 4.315 0.930 ;
        RECT  4.220 2.135 4.225 2.295 ;
        RECT  4.060 1.980 4.220 2.295 ;
        RECT  3.220 0.770 4.155 0.930 ;
        RECT  3.560 1.980 4.060 2.140 ;
        RECT  3.745 1.450 4.005 1.710 ;
        RECT  3.540 1.110 3.560 2.140 ;
        RECT  3.400 1.110 3.540 2.190 ;
        RECT  3.380 2.370 3.540 2.735 ;
        RECT  3.380 1.930 3.400 2.190 ;
        RECT  3.195 2.370 3.380 2.530 ;
        RECT  3.195 0.770 3.220 1.595 ;
        RECT  3.060 0.770 3.195 2.530 ;
        RECT  3.005 3.100 3.140 3.260 ;
        RECT  3.035 1.350 3.060 2.530 ;
        RECT  2.850 2.730 3.005 3.260 ;
        RECT  2.850 0.925 2.880 1.185 ;
        RECT  2.845 0.925 2.850 3.260 ;
        RECT  2.690 0.925 2.845 2.890 ;
        RECT  2.370 0.870 2.510 2.920 ;
        RECT  2.350 0.585 2.370 2.920 ;
        RECT  2.210 0.585 2.350 1.125 ;
        RECT  2.225 2.320 2.350 2.920 ;
        RECT  0.825 2.760 2.225 2.920 ;
        RECT  0.605 0.585 2.210 0.745 ;
        RECT  2.030 1.410 2.170 1.670 ;
        RECT  1.870 0.925 2.030 1.670 ;
        RECT  0.970 0.925 1.870 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.665 0.925 0.825 2.215 ;
        RECT  0.565 2.645 0.825 2.920 ;
        RECT  0.445 0.455 0.605 0.745 ;
    END
END SDFFSRX2

MACRO SDFFSRX1
    CLASS CORE ;
    FOREIGN SDFFSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.910 2.520 9.995 2.810 ;
        RECT  9.785 2.520 9.910 3.260 ;
        RECT  9.750 2.585 9.785 3.260 ;
        RECT  9.630 3.000 9.750 3.260 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.010 1.600 1.320 2.020 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.1105 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.805 5.865 2.065 ;
        RECT  5.495 1.700 5.855 2.065 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.370 2.335 11.375 2.810 ;
        RECT  11.210 0.645 11.370 2.810 ;
        RECT  11.165 0.645 11.210 0.945 ;
        RECT  11.165 2.335 11.210 2.810 ;
        RECT  10.905 0.645 11.165 0.805 ;
        RECT  10.920 2.595 11.165 2.810 ;
        RECT  10.660 2.595 10.920 3.195 ;
        RECT  10.645 0.545 10.905 0.805 ;
        END
        ANTENNADIFFAREA     0.3838 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.625 0.920 11.835 2.750 ;
        RECT  11.575 0.920 11.625 1.180 ;
        RECT  11.575 2.150 11.625 2.750 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.675 1.925 1.715 2.500 ;
        RECT  1.515 1.265 1.675 2.500 ;
        RECT  1.390 1.265 1.515 1.425 ;
        RECT  1.505 1.925 1.515 2.500 ;
        RECT  1.235 2.240 1.505 2.500 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 1.695 4.935 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.435 -0.250 11.960 0.250 ;
        RECT  11.175 -0.250 11.435 0.405 ;
        RECT  10.355 -0.250 11.175 0.250 ;
        RECT  10.095 -0.250 10.355 0.405 ;
        RECT  5.600 -0.250 10.095 0.250 ;
        RECT  5.340 -0.250 5.600 0.405 ;
        RECT  3.870 -0.250 5.340 0.250 ;
        RECT  3.610 -0.250 3.870 0.405 ;
        RECT  1.550 -0.250 3.610 0.250 ;
        RECT  1.290 -0.250 1.550 0.405 ;
        RECT  0.270 -0.250 1.290 0.250 ;
        RECT  0.270 1.035 0.335 1.295 ;
        RECT  0.110 -0.250 0.270 1.295 ;
        RECT  0.000 -0.250 0.110 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.435 3.440 11.960 3.940 ;
        RECT  11.175 3.285 11.435 3.940 ;
        RECT  10.355 3.440 11.175 3.940 ;
        RECT  10.175 2.765 10.355 3.940 ;
        RECT  10.095 3.285 10.175 3.940 ;
        RECT  8.085 3.440 10.095 3.940 ;
        RECT  7.825 3.285 8.085 3.940 ;
        RECT  6.345 3.440 7.825 3.940 ;
        RECT  5.405 3.055 6.345 3.940 ;
        RECT  3.840 3.440 5.405 3.940 ;
        RECT  3.580 2.900 3.840 3.940 ;
        RECT  1.555 3.440 3.580 3.940 ;
        RECT  1.295 3.285 1.555 3.940 ;
        RECT  0.385 3.440 1.295 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.940 1.635 11.030 1.895 ;
        RECT  10.780 1.120 10.940 2.345 ;
        RECT  10.715 1.120 10.780 1.380 ;
        RECT  10.665 1.900 10.780 2.345 ;
        RECT  9.580 1.900 10.665 2.060 ;
        RECT  10.500 1.560 10.600 1.720 ;
        RECT  10.340 1.275 10.500 1.720 ;
        RECT  8.890 1.275 10.340 1.435 ;
        RECT  9.850 0.835 9.950 1.095 ;
        RECT  9.690 0.475 9.850 1.095 ;
        RECT  7.280 0.475 9.690 0.635 ;
        RECT  9.420 1.615 9.580 2.060 ;
        RECT  9.195 2.255 9.455 2.515 ;
        RECT  9.320 1.615 9.420 1.875 ;
        RECT  9.060 0.815 9.220 1.095 ;
        RECT  9.150 2.355 9.195 2.515 ;
        RECT  8.990 2.355 9.150 3.100 ;
        RECT  8.130 0.815 9.060 0.975 ;
        RECT  6.990 2.940 8.990 3.100 ;
        RECT  8.810 1.615 8.910 1.775 ;
        RECT  8.615 1.175 8.890 1.435 ;
        RECT  8.650 1.615 8.810 2.755 ;
        RECT  6.600 2.595 8.650 2.755 ;
        RECT  8.470 1.275 8.615 1.435 ;
        RECT  8.310 1.275 8.470 2.340 ;
        RECT  8.165 2.080 8.310 2.340 ;
        RECT  7.985 0.815 8.130 1.655 ;
        RECT  7.970 0.815 7.985 1.935 ;
        RECT  7.885 1.495 7.970 1.935 ;
        RECT  7.825 1.495 7.885 2.410 ;
        RECT  7.725 1.675 7.825 2.410 ;
        RECT  7.630 0.815 7.790 1.285 ;
        RECT  6.945 2.250 7.725 2.410 ;
        RECT  7.385 1.125 7.630 1.285 ;
        RECT  7.225 1.125 7.385 2.050 ;
        RECT  7.120 0.475 7.280 0.945 ;
        RECT  6.940 1.125 7.225 1.285 ;
        RECT  7.125 1.790 7.225 2.050 ;
        RECT  6.830 2.940 6.990 3.210 ;
        RECT  6.785 1.465 6.945 2.410 ;
        RECT  6.780 0.590 6.940 1.285 ;
        RECT  6.675 3.050 6.830 3.210 ;
        RECT  6.600 1.465 6.785 1.625 ;
        RECT  4.935 0.590 6.780 0.750 ;
        RECT  6.440 0.930 6.600 1.625 ;
        RECT  6.260 1.860 6.600 2.120 ;
        RECT  6.440 2.595 6.600 2.870 ;
        RECT  5.275 0.930 6.440 1.090 ;
        RECT  4.520 2.710 6.440 2.870 ;
        RECT  6.100 1.270 6.260 2.425 ;
        RECT  5.770 1.270 6.100 1.430 ;
        RECT  5.730 2.265 6.100 2.425 ;
        RECT  5.115 0.930 5.275 2.355 ;
        RECT  4.250 1.270 5.115 1.430 ;
        RECT  4.715 2.195 5.115 2.355 ;
        RECT  4.825 3.050 5.085 3.260 ;
        RECT  4.775 0.590 4.935 1.090 ;
        RECT  4.180 3.050 4.825 3.210 ;
        RECT  3.765 0.930 4.775 1.090 ;
        RECT  4.360 2.215 4.520 2.870 ;
        RECT  4.200 0.490 4.460 0.750 ;
        RECT  3.585 2.215 4.360 2.375 ;
        RECT  4.090 1.270 4.250 2.035 ;
        RECT  3.325 0.590 4.200 0.750 ;
        RECT  4.020 2.560 4.180 3.210 ;
        RECT  3.990 1.775 4.090 2.035 ;
        RECT  3.160 2.560 4.020 2.720 ;
        RECT  3.605 0.930 3.765 1.455 ;
        RECT  3.505 1.195 3.605 1.455 ;
        RECT  3.425 2.100 3.585 2.375 ;
        RECT  3.100 2.100 3.425 2.260 ;
        RECT  3.165 0.590 3.325 1.420 ;
        RECT  3.100 1.260 3.165 1.420 ;
        RECT  2.900 2.440 3.160 2.720 ;
        RECT  2.940 1.260 3.100 2.260 ;
        RECT  2.760 0.820 2.975 1.080 ;
        RECT  2.760 2.440 2.900 2.600 ;
        RECT  2.715 0.820 2.760 2.600 ;
        RECT  2.600 0.920 2.715 2.600 ;
        RECT  2.420 2.780 2.485 3.040 ;
        RECT  2.260 0.585 2.420 3.040 ;
        RECT  2.195 0.585 2.260 1.085 ;
        RECT  2.225 2.715 2.260 3.040 ;
        RECT  0.845 2.715 2.225 2.875 ;
        RECT  0.610 0.585 2.195 0.745 ;
        RECT  2.015 1.265 2.080 1.525 ;
        RECT  1.855 0.925 2.015 1.525 ;
        RECT  0.970 0.925 1.855 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.585 2.615 0.845 2.875 ;
        RECT  0.665 0.925 0.825 2.285 ;
        RECT  0.450 0.440 0.610 0.745 ;
    END
END SDFFSRX1

MACRO SDFFSRXL
    CLASS CORE ;
    FOREIGN SDFFSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.910 2.520 9.995 2.810 ;
        RECT  9.785 2.520 9.910 3.260 ;
        RECT  9.750 2.585 9.785 3.260 ;
        RECT  9.630 3.000 9.750 3.260 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.010 1.600 1.320 2.020 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.530 1.655 5.855 2.065 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.370 2.335 11.375 2.810 ;
        RECT  11.210 0.710 11.370 2.810 ;
        RECT  11.165 0.710 11.210 0.945 ;
        RECT  11.165 2.335 11.210 2.810 ;
        RECT  10.930 0.710 11.165 0.870 ;
        RECT  10.630 2.550 11.165 2.810 ;
        RECT  10.670 0.610 10.930 0.870 ;
        END
        ANTENNADIFFAREA     0.2135 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.810 0.695 11.835 2.570 ;
        RECT  11.625 0.535 11.810 2.570 ;
        RECT  11.550 0.535 11.625 0.795 ;
        RECT  11.575 2.310 11.625 2.570 ;
        END
        ANTENNADIFFAREA     0.2898 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.250 1.720 2.510 ;
        RECT  1.675 1.925 1.715 2.510 ;
        RECT  1.515 1.265 1.675 2.510 ;
        RECT  1.390 1.265 1.515 1.425 ;
        RECT  1.505 1.925 1.515 2.510 ;
        RECT  1.235 2.250 1.505 2.510 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 1.695 4.935 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.350 -0.250 11.960 0.250 ;
        RECT  10.090 -0.250 10.350 0.405 ;
        RECT  5.600 -0.250 10.090 0.250 ;
        RECT  5.340 -0.250 5.600 0.405 ;
        RECT  3.825 -0.250 5.340 0.250 ;
        RECT  3.565 -0.250 3.825 0.405 ;
        RECT  1.550 -0.250 3.565 0.250 ;
        RECT  1.290 -0.250 1.550 0.405 ;
        RECT  0.265 -0.250 1.290 0.250 ;
        RECT  0.265 1.035 0.335 1.295 ;
        RECT  0.105 -0.250 0.265 1.295 ;
        RECT  0.000 -0.250 0.105 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.435 3.440 11.960 3.940 ;
        RECT  11.175 3.285 11.435 3.940 ;
        RECT  10.350 3.440 11.175 3.940 ;
        RECT  10.090 3.285 10.350 3.940 ;
        RECT  8.085 3.440 10.090 3.940 ;
        RECT  7.825 3.285 8.085 3.940 ;
        RECT  6.345 3.440 7.825 3.940 ;
        RECT  5.405 3.055 6.345 3.940 ;
        RECT  3.890 3.440 5.405 3.940 ;
        RECT  3.630 2.900 3.890 3.940 ;
        RECT  1.555 3.440 3.630 3.940 ;
        RECT  1.295 3.285 1.555 3.940 ;
        RECT  0.385 3.440 1.295 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.940 1.635 11.030 1.895 ;
        RECT  10.920 1.120 10.940 2.085 ;
        RECT  10.780 1.120 10.920 2.300 ;
        RECT  10.720 1.120 10.780 1.380 ;
        RECT  10.660 1.920 10.780 2.300 ;
        RECT  9.580 1.920 10.660 2.080 ;
        RECT  10.500 1.560 10.600 1.720 ;
        RECT  10.340 1.275 10.500 1.720 ;
        RECT  8.890 1.275 10.340 1.435 ;
        RECT  9.850 0.835 9.950 1.095 ;
        RECT  9.690 0.475 9.850 1.095 ;
        RECT  7.220 0.475 9.690 0.635 ;
        RECT  9.320 1.820 9.580 2.080 ;
        RECT  9.195 2.265 9.455 2.525 ;
        RECT  9.060 0.835 9.220 1.095 ;
        RECT  9.150 2.365 9.195 2.525 ;
        RECT  8.990 2.365 9.150 3.100 ;
        RECT  8.130 0.835 9.060 0.995 ;
        RECT  6.980 2.940 8.990 3.100 ;
        RECT  8.810 1.615 8.940 1.775 ;
        RECT  8.615 1.175 8.890 1.435 ;
        RECT  8.650 1.615 8.810 2.755 ;
        RECT  6.600 2.595 8.650 2.755 ;
        RECT  8.470 1.275 8.615 1.435 ;
        RECT  8.310 1.275 8.470 2.395 ;
        RECT  8.130 2.135 8.310 2.395 ;
        RECT  7.970 0.835 8.130 1.910 ;
        RECT  7.950 1.750 7.970 1.910 ;
        RECT  7.850 1.750 7.950 2.050 ;
        RECT  7.690 1.750 7.850 2.410 ;
        RECT  7.630 0.870 7.790 1.480 ;
        RECT  6.940 2.250 7.690 2.410 ;
        RECT  7.380 1.320 7.630 1.480 ;
        RECT  7.220 1.320 7.380 2.050 ;
        RECT  7.060 0.475 7.220 1.130 ;
        RECT  6.880 1.320 7.220 1.480 ;
        RECT  7.120 1.790 7.220 2.050 ;
        RECT  6.780 2.940 6.980 3.210 ;
        RECT  6.780 1.660 6.940 2.410 ;
        RECT  6.720 0.590 6.880 1.480 ;
        RECT  6.540 1.660 6.780 1.820 ;
        RECT  6.720 3.050 6.780 3.210 ;
        RECT  4.935 0.590 6.720 0.750 ;
        RECT  6.200 2.000 6.600 2.260 ;
        RECT  6.440 2.595 6.600 2.870 ;
        RECT  6.380 0.930 6.540 1.820 ;
        RECT  4.570 2.710 6.440 2.870 ;
        RECT  5.275 0.930 6.380 1.090 ;
        RECT  6.040 1.270 6.200 2.425 ;
        RECT  5.770 1.270 6.040 1.430 ;
        RECT  5.770 2.265 6.040 2.425 ;
        RECT  5.115 0.930 5.275 2.355 ;
        RECT  4.250 1.270 5.115 1.430 ;
        RECT  4.755 2.195 5.115 2.355 ;
        RECT  4.825 3.050 5.085 3.255 ;
        RECT  4.775 0.590 4.935 1.090 ;
        RECT  4.230 3.050 4.825 3.210 ;
        RECT  3.765 0.930 4.775 1.090 ;
        RECT  4.410 2.215 4.570 2.870 ;
        RECT  4.200 0.490 4.460 0.750 ;
        RECT  3.635 2.215 4.410 2.375 ;
        RECT  4.090 1.270 4.250 2.035 ;
        RECT  4.070 2.560 4.230 3.210 ;
        RECT  3.325 0.590 4.200 0.750 ;
        RECT  3.990 1.775 4.090 2.035 ;
        RECT  3.160 2.560 4.070 2.720 ;
        RECT  3.605 0.930 3.765 1.455 ;
        RECT  3.475 2.100 3.635 2.375 ;
        RECT  3.505 1.195 3.605 1.455 ;
        RECT  3.100 2.100 3.475 2.260 ;
        RECT  3.165 0.590 3.325 1.420 ;
        RECT  3.100 1.260 3.165 1.420 ;
        RECT  2.900 2.440 3.160 2.720 ;
        RECT  2.940 1.260 3.100 2.260 ;
        RECT  2.760 0.820 2.975 1.080 ;
        RECT  2.760 2.440 2.900 2.600 ;
        RECT  2.715 0.820 2.760 2.600 ;
        RECT  2.600 0.920 2.715 2.600 ;
        RECT  2.420 2.780 2.485 3.040 ;
        RECT  2.260 0.585 2.420 3.040 ;
        RECT  2.195 0.585 2.260 1.085 ;
        RECT  2.225 2.720 2.260 3.040 ;
        RECT  0.810 2.720 2.225 2.880 ;
        RECT  0.605 0.585 2.195 0.745 ;
        RECT  2.015 1.265 2.080 1.525 ;
        RECT  1.855 0.925 2.015 1.525 ;
        RECT  0.970 0.925 1.855 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.665 0.925 0.825 2.285 ;
        RECT  0.550 2.620 0.810 2.880 ;
        RECT  0.445 0.440 0.605 0.745 ;
    END
END SDFFSRXL

MACRO SDFFSX4
    CLASS CORE ;
    FOREIGN SDFFSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.340 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.325 2.020 9.585 2.400 ;
        RECT  8.945 2.240 9.325 2.400 ;
        RECT  8.785 2.240 8.945 3.260 ;
        RECT  8.535 3.100 8.785 3.260 ;
        END
        ANTENNAGATEAREA     0.3302 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.545 1.295 1.990 ;
        END
        ANTENNAGATEAREA     0.0793 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.1716 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.380 0.695 11.480 1.295 ;
        RECT  11.215 0.695 11.380 2.555 ;
        RECT  11.165 0.695 11.215 1.580 ;
        END
        ANTENNADIFFAREA     0.7543 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.660 1.105 12.755 2.585 ;
        RECT  12.400 0.595 12.660 2.750 ;
        END
        ANTENNADIFFAREA     0.7258 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.265 1.735 1.425 ;
        RECT  1.475 1.265 1.715 2.425 ;
        RECT  1.215 2.170 1.475 2.425 ;
        END
        ANTENNAGATEAREA     0.1560 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.700 4.395 2.240 ;
        END
        ANTENNAGATEAREA     0.0650 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.210 -0.250 13.340 0.250 ;
        RECT  12.950 -0.250 13.210 1.195 ;
        RECT  12.110 -0.250 12.950 0.250 ;
        RECT  11.850 -0.250 12.110 1.195 ;
        RECT  10.980 -0.250 11.850 0.250 ;
        RECT  10.720 -0.250 10.980 1.195 ;
        RECT  9.415 -0.250 10.720 0.250 ;
        RECT  9.155 -0.250 9.415 1.075 ;
        RECT  6.760 -0.250 9.155 0.250 ;
        RECT  6.500 -0.250 6.760 0.405 ;
        RECT  4.045 -0.250 6.500 0.250 ;
        RECT  3.785 -0.250 4.045 0.405 ;
        RECT  1.605 -0.250 3.785 0.250 ;
        RECT  1.345 -0.250 1.605 0.405 ;
        RECT  0.285 -0.250 1.345 0.250 ;
        RECT  0.285 1.035 0.385 1.295 ;
        RECT  0.125 -0.250 0.285 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.210 3.440 13.340 3.940 ;
        RECT  12.950 2.120 13.210 3.940 ;
        RECT  12.110 3.440 12.950 3.940 ;
        RECT  11.900 2.155 12.110 3.940 ;
        RECT  11.850 3.285 11.900 3.940 ;
        RECT  10.795 3.440 11.850 3.940 ;
        RECT  10.695 3.285 10.795 3.940 ;
        RECT  10.535 2.240 10.695 3.940 ;
        RECT  9.445 3.440 10.535 3.940 ;
        RECT  9.445 2.585 9.625 2.845 ;
        RECT  9.185 2.585 9.445 3.940 ;
        RECT  7.795 3.440 9.185 3.940 ;
        RECT  7.535 3.285 7.795 3.940 ;
        RECT  5.640 3.440 7.535 3.940 ;
        RECT  5.040 3.105 5.640 3.940 ;
        RECT  4.145 3.440 5.040 3.940 ;
        RECT  3.885 3.105 4.145 3.940 ;
        RECT  1.745 3.440 3.885 3.940 ;
        RECT  1.485 3.285 1.745 3.940 ;
        RECT  0.385 3.440 1.485 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.055 1.520 12.215 1.925 ;
        RECT  11.720 1.765 12.055 1.925 ;
        RECT  11.560 1.765 11.720 2.915 ;
        RECT  11.035 2.755 11.560 2.915 ;
        RECT  10.875 1.885 11.035 2.915 ;
        RECT  10.355 1.885 10.875 2.045 ;
        RECT  10.355 0.965 10.440 1.225 ;
        RECT  10.235 0.965 10.355 2.400 ;
        RECT  10.195 0.965 10.235 2.840 ;
        RECT  10.180 0.965 10.195 1.225 ;
        RECT  10.135 2.240 10.195 2.840 ;
        RECT  9.975 2.240 10.135 3.190 ;
        RECT  9.855 1.675 10.015 1.960 ;
        RECT  9.625 3.030 9.975 3.190 ;
        RECT  9.665 0.555 9.925 1.495 ;
        RECT  8.475 1.675 9.855 1.835 ;
        RECT  8.905 1.335 9.665 1.495 ;
        RECT  8.855 0.555 8.905 1.495 ;
        RECT  8.665 0.480 8.855 1.495 ;
        RECT  7.100 0.480 8.665 0.640 ;
        RECT  8.315 0.910 8.475 2.920 ;
        RECT  7.885 0.910 8.315 1.085 ;
        RECT  8.200 2.660 8.315 2.920 ;
        RECT  7.755 2.660 8.200 2.820 ;
        RECT  7.975 1.830 8.135 2.475 ;
        RECT  7.465 1.830 7.975 1.990 ;
        RECT  7.625 0.825 7.885 1.085 ;
        RECT  7.595 2.175 7.755 3.100 ;
        RECT  6.475 2.940 7.595 3.100 ;
        RECT  7.445 1.425 7.465 1.990 ;
        RECT  7.415 1.270 7.445 1.990 ;
        RECT  7.255 1.270 7.415 2.760 ;
        RECT  6.115 0.925 7.315 1.085 ;
        RECT  7.205 1.270 7.255 1.685 ;
        RECT  6.275 2.600 7.255 2.760 ;
        RECT  6.545 1.270 7.205 1.430 ;
        RECT  6.940 0.480 7.100 0.745 ;
        RECT  6.975 2.255 7.075 2.415 ;
        RECT  6.815 1.620 6.975 2.415 ;
        RECT  6.305 0.585 6.940 0.745 ;
        RECT  6.115 1.620 6.815 1.780 ;
        RECT  5.590 1.970 6.625 2.130 ;
        RECT  6.315 2.940 6.475 3.215 ;
        RECT  6.145 0.470 6.305 0.745 ;
        RECT  6.130 2.380 6.275 2.760 ;
        RECT  5.575 0.470 6.145 0.630 ;
        RECT  5.970 2.380 6.130 3.260 ;
        RECT  5.825 0.925 6.115 1.780 ;
        RECT  5.825 3.050 5.970 3.260 ;
        RECT  5.135 1.620 5.825 1.780 ;
        RECT  5.430 1.970 5.590 2.920 ;
        RECT  5.315 0.470 5.575 1.100 ;
        RECT  3.605 2.760 5.430 2.920 ;
        RECT  5.115 1.980 5.145 2.580 ;
        RECT  5.115 1.015 5.135 1.780 ;
        RECT  4.955 1.015 5.115 2.580 ;
        RECT  4.805 1.015 4.955 1.280 ;
        RECT  3.915 1.120 4.805 1.280 ;
        RECT  4.615 1.495 4.775 2.580 ;
        RECT  4.365 0.545 4.625 0.745 ;
        RECT  3.285 2.420 4.615 2.580 ;
        RECT  2.980 0.585 4.365 0.745 ;
        RECT  3.705 1.120 3.915 1.515 ;
        RECT  3.655 1.255 3.705 1.515 ;
        RECT  3.345 2.760 3.605 3.020 ;
        RECT  2.945 2.760 3.345 2.920 ;
        RECT  3.125 0.925 3.285 2.580 ;
        RECT  3.025 0.925 3.125 1.185 ;
        RECT  2.845 0.495 2.980 0.745 ;
        RECT  2.845 1.485 2.945 2.920 ;
        RECT  2.785 0.495 2.845 2.920 ;
        RECT  2.685 0.495 2.785 1.645 ;
        RECT  2.505 1.930 2.605 2.885 ;
        RECT  2.445 0.585 2.505 2.885 ;
        RECT  2.345 0.585 2.445 2.090 ;
        RECT  0.785 2.725 2.445 2.885 ;
        RECT  0.725 0.585 2.345 0.745 ;
        RECT  2.005 0.925 2.165 1.635 ;
        RECT  0.970 0.925 2.005 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.665 0.925 0.825 2.215 ;
        RECT  0.525 2.725 0.785 2.985 ;
        RECT  0.465 0.430 0.725 0.745 ;
    END
END SDFFSX4

MACRO SDFFSX2
    CLASS CORE ;
    FOREIGN SDFFSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.685 2.160 8.945 2.420 ;
        RECT  8.615 2.160 8.685 2.400 ;
        RECT  8.405 2.110 8.615 2.400 ;
        RECT  8.175 2.240 8.405 2.400 ;
        RECT  8.015 2.240 8.175 3.185 ;
        RECT  7.665 3.025 8.015 3.185 ;
        RECT  7.400 3.025 7.665 3.255 ;
        END
        ANTENNAGATEAREA     0.1898 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.595 1.295 2.045 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.085 0.695 10.245 1.295 ;
        RECT  9.780 0.695 10.085 2.555 ;
        END
        ANTENNADIFFAREA     0.7460 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.115 0.595 11.375 3.045 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.270 1.735 1.530 ;
        RECT  1.545 1.270 1.715 2.400 ;
        RECT  1.505 1.270 1.545 2.535 ;
        RECT  1.475 1.270 1.505 1.530 ;
        RECT  1.285 2.240 1.505 2.535 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.740 4.250 2.035 ;
        RECT  3.805 1.700 4.015 2.035 ;
        RECT  3.765 1.740 3.805 2.035 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.825 -0.250 11.500 0.250 ;
        RECT  10.565 -0.250 10.825 1.195 ;
        RECT  8.945 -0.250 10.565 0.250 ;
        RECT  8.685 -0.250 8.945 1.435 ;
        RECT  5.275 -0.250 8.685 0.250 ;
        RECT  5.015 -0.250 5.275 0.405 ;
        RECT  4.045 -0.250 5.015 0.250 ;
        RECT  3.785 -0.250 4.045 0.405 ;
        RECT  1.605 -0.250 3.785 0.250 ;
        RECT  1.345 -0.250 1.605 0.405 ;
        RECT  0.280 -0.250 1.345 0.250 ;
        RECT  0.280 1.035 0.385 1.295 ;
        RECT  0.120 -0.250 0.280 1.295 ;
        RECT  0.000 -0.250 0.120 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.825 3.440 11.500 3.940 ;
        RECT  10.615 2.120 10.825 3.940 ;
        RECT  10.565 3.285 10.615 3.940 ;
        RECT  8.985 3.440 10.565 3.940 ;
        RECT  8.725 2.945 8.985 3.940 ;
        RECT  7.220 3.440 8.725 3.940 ;
        RECT  6.960 3.035 7.220 3.940 ;
        RECT  5.310 3.440 6.960 3.940 ;
        RECT  5.050 3.105 5.310 3.940 ;
        RECT  4.045 3.440 5.050 3.940 ;
        RECT  3.785 3.105 4.045 3.940 ;
        RECT  1.745 3.440 3.785 3.940 ;
        RECT  1.485 3.285 1.745 3.940 ;
        RECT  0.385 3.440 1.485 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.770 1.520 10.930 1.810 ;
        RECT  10.435 1.650 10.770 1.810 ;
        RECT  10.275 1.650 10.435 3.025 ;
        RECT  9.595 2.865 10.275 3.025 ;
        RECT  9.545 2.765 9.595 3.025 ;
        RECT  9.385 1.035 9.545 3.025 ;
        RECT  9.255 1.035 9.385 1.295 ;
        RECT  9.335 2.605 9.385 3.025 ;
        RECT  8.515 2.605 9.335 2.765 ;
        RECT  9.045 1.680 9.205 1.940 ;
        RECT  7.835 1.680 9.045 1.840 ;
        RECT  8.355 2.605 8.515 3.260 ;
        RECT  8.175 0.470 8.435 1.435 ;
        RECT  5.620 0.470 8.175 0.630 ;
        RECT  7.675 0.915 7.835 2.845 ;
        RECT  7.485 0.915 7.675 1.075 ;
        RECT  7.125 2.685 7.675 2.845 ;
        RECT  7.335 1.355 7.495 2.340 ;
        RECT  7.225 0.815 7.485 1.075 ;
        RECT  7.115 1.355 7.335 1.515 ;
        RECT  6.965 2.085 7.125 2.845 ;
        RECT  6.855 1.255 7.115 1.515 ;
        RECT  6.655 0.815 6.915 1.075 ;
        RECT  6.775 1.355 6.855 1.515 ;
        RECT  6.615 1.355 6.775 3.220 ;
        RECT  6.010 0.815 6.655 0.980 ;
        RECT  6.355 1.355 6.615 1.515 ;
        RECT  5.990 3.060 6.615 3.220 ;
        RECT  6.275 1.695 6.435 2.845 ;
        RECT  6.195 1.160 6.355 1.515 ;
        RECT  6.010 1.695 6.275 1.855 ;
        RECT  5.470 2.040 6.020 2.200 ;
        RECT  5.850 0.815 6.010 1.855 ;
        RECT  5.830 3.000 5.990 3.260 ;
        RECT  5.585 1.015 5.850 1.275 ;
        RECT  5.670 2.510 5.830 3.260 ;
        RECT  5.460 0.470 5.620 0.815 ;
        RECT  5.425 1.015 5.585 1.505 ;
        RECT  5.310 2.040 5.470 2.920 ;
        RECT  5.175 0.655 5.460 0.815 ;
        RECT  4.615 1.345 5.425 1.505 ;
        RECT  4.615 2.760 5.310 2.920 ;
        RECT  5.015 0.655 5.175 1.165 ;
        RECT  5.105 1.690 5.110 1.850 ;
        RECT  4.945 1.690 5.105 2.580 ;
        RECT  4.915 0.905 5.015 1.165 ;
        RECT  4.850 1.690 4.945 1.850 ;
        RECT  3.185 2.420 4.945 2.580 ;
        RECT  4.615 2.080 4.740 2.240 ;
        RECT  4.365 0.445 4.625 0.745 ;
        RECT  4.455 1.015 4.615 2.240 ;
        RECT  4.355 2.760 4.615 3.020 ;
        RECT  3.655 1.345 4.455 1.505 ;
        RECT  2.845 0.585 4.365 0.745 ;
        RECT  3.460 2.760 4.355 2.920 ;
        RECT  3.200 2.760 3.460 3.025 ;
        RECT  2.845 2.760 3.200 2.920 ;
        RECT  3.025 0.925 3.185 2.580 ;
        RECT  2.685 0.585 2.845 2.920 ;
        RECT  2.345 0.535 2.505 3.105 ;
        RECT  0.720 0.585 2.345 0.745 ;
        RECT  0.895 2.945 2.345 3.105 ;
        RECT  2.005 0.925 2.165 1.715 ;
        RECT  0.970 0.925 2.005 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.635 2.725 0.895 3.105 ;
        RECT  0.665 0.925 0.825 2.305 ;
        RECT  0.460 0.430 0.720 0.745 ;
    END
END SDFFSX2

MACRO SDFFSX1
    CLASS CORE ;
    FOREIGN SDFFSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.405 1.515 8.615 1.990 ;
        RECT  8.345 1.515 8.405 1.775 ;
        RECT  8.175 1.615 8.345 1.775 ;
        RECT  8.015 1.615 8.175 3.205 ;
        RECT  7.665 3.045 8.015 3.205 ;
        RECT  7.405 3.045 7.665 3.255 ;
        END
        ANTENNAGATEAREA     0.1144 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.595 1.295 2.045 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.995 0.655 10.010 2.755 ;
        RECT  9.850 0.655 9.995 2.810 ;
        RECT  9.475 0.655 9.850 0.815 ;
        RECT  9.785 2.520 9.850 2.810 ;
        RECT  9.545 2.595 9.785 2.810 ;
        RECT  9.285 2.595 9.545 3.195 ;
        RECT  9.215 0.555 9.475 0.815 ;
        END
        ANTENNADIFFAREA     0.3796 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.195 0.975 10.455 2.750 ;
        END
        ANTENNADIFFAREA     0.3772 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.270 1.735 1.530 ;
        RECT  1.505 1.270 1.715 2.435 ;
        RECT  1.475 1.270 1.505 1.530 ;
        RECT  1.475 2.275 1.505 2.435 ;
        RECT  1.215 2.275 1.475 2.535 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.740 4.250 2.035 ;
        RECT  3.805 1.700 4.015 2.035 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.015 -0.250 10.580 0.250 ;
        RECT  9.755 -0.250 10.015 0.405 ;
        RECT  8.935 -0.250 9.755 0.250 ;
        RECT  8.675 -0.250 8.935 0.795 ;
        RECT  5.245 -0.250 8.675 0.250 ;
        RECT  4.985 -0.250 5.245 0.405 ;
        RECT  4.045 -0.250 4.985 0.250 ;
        RECT  3.785 -0.250 4.045 0.405 ;
        RECT  1.540 -0.250 3.785 0.250 ;
        RECT  1.280 -0.250 1.540 0.405 ;
        RECT  0.265 -0.250 1.280 0.250 ;
        RECT  0.265 1.035 0.385 1.295 ;
        RECT  0.105 -0.250 0.265 1.295 ;
        RECT  0.000 -0.250 0.105 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.055 3.440 10.580 3.940 ;
        RECT  9.795 3.285 10.055 3.940 ;
        RECT  8.975 3.440 9.795 3.940 ;
        RECT  8.715 2.735 8.975 3.940 ;
        RECT  7.220 3.440 8.715 3.940 ;
        RECT  6.960 2.985 7.220 3.940 ;
        RECT  5.310 3.440 6.960 3.940 ;
        RECT  5.050 3.105 5.310 3.940 ;
        RECT  4.045 3.440 5.050 3.940 ;
        RECT  3.785 3.105 4.045 3.940 ;
        RECT  1.675 3.440 3.785 3.940 ;
        RECT  1.415 3.285 1.675 3.940 ;
        RECT  0.385 3.440 1.415 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.545 1.125 9.670 2.245 ;
        RECT  9.510 1.125 9.545 2.345 ;
        RECT  9.295 1.125 9.510 1.385 ;
        RECT  9.285 2.085 9.510 2.345 ;
        RECT  8.615 2.185 9.285 2.345 ;
        RECT  9.055 1.560 9.155 1.820 ;
        RECT  8.895 1.170 9.055 1.820 ;
        RECT  7.835 1.170 8.895 1.330 ;
        RECT  8.355 2.180 8.615 2.440 ;
        RECT  8.225 0.730 8.325 0.990 ;
        RECT  8.065 0.470 8.225 0.990 ;
        RECT  5.585 0.470 8.065 0.630 ;
        RECT  7.675 0.910 7.835 2.835 ;
        RECT  7.185 0.910 7.675 1.070 ;
        RECT  7.550 2.575 7.675 2.835 ;
        RECT  7.125 2.575 7.550 2.735 ;
        RECT  7.335 1.280 7.495 2.395 ;
        RECT  6.775 1.280 7.335 1.440 ;
        RECT  6.965 2.085 7.125 2.735 ;
        RECT  6.615 0.810 6.875 1.100 ;
        RECT  6.615 1.280 6.775 3.220 ;
        RECT  5.925 0.810 6.615 0.970 ;
        RECT  6.365 1.280 6.615 1.440 ;
        RECT  5.880 3.060 6.615 3.220 ;
        RECT  6.275 1.620 6.435 2.845 ;
        RECT  6.105 1.150 6.365 1.440 ;
        RECT  5.925 1.620 6.275 1.780 ;
        RECT  5.280 1.960 6.020 2.120 ;
        RECT  5.765 0.810 5.925 1.780 ;
        RECT  5.750 2.300 5.880 3.220 ;
        RECT  4.665 1.345 5.765 1.505 ;
        RECT  5.620 2.300 5.750 3.260 ;
        RECT  5.490 3.000 5.620 3.260 ;
        RECT  5.425 0.470 5.585 1.065 ;
        RECT  5.255 0.905 5.425 1.065 ;
        RECT  5.120 1.960 5.280 2.890 ;
        RECT  4.995 0.905 5.255 1.165 ;
        RECT  4.615 2.730 5.120 2.890 ;
        RECT  3.185 2.390 4.940 2.550 ;
        RECT  4.615 2.005 4.740 2.165 ;
        RECT  4.615 1.015 4.665 1.505 ;
        RECT  4.365 0.445 4.625 0.745 ;
        RECT  4.455 1.015 4.615 2.165 ;
        RECT  4.355 2.730 4.615 2.990 ;
        RECT  4.405 1.015 4.455 1.505 ;
        RECT  3.655 1.345 4.405 1.505 ;
        RECT  2.845 0.585 4.365 0.745 ;
        RECT  3.435 2.730 4.355 2.890 ;
        RECT  3.175 2.730 3.435 2.990 ;
        RECT  3.025 0.925 3.185 2.550 ;
        RECT  2.845 2.730 3.175 2.890 ;
        RECT  2.685 0.585 2.845 2.890 ;
        RECT  2.345 0.430 2.505 2.875 ;
        RECT  0.605 0.585 2.345 0.745 ;
        RECT  0.795 2.715 2.345 2.875 ;
        RECT  2.005 0.925 2.165 1.530 ;
        RECT  0.970 0.925 2.005 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.665 0.925 0.825 2.305 ;
        RECT  0.535 2.660 0.795 2.920 ;
        RECT  0.445 0.430 0.605 0.745 ;
    END
END SDFFSX1

MACRO SDFFSXL
    CLASS CORE ;
    FOREIGN SDFFSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.345 1.515 8.615 1.990 ;
        RECT  8.175 1.830 8.345 1.990 ;
        RECT  8.015 1.830 8.175 3.255 ;
        RECT  7.405 3.095 8.015 3.255 ;
        END
        ANTENNAGATEAREA     0.0793 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.595 1.295 2.045 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.850 0.710 10.010 2.810 ;
        RECT  9.510 0.710 9.850 0.870 ;
        RECT  9.785 2.520 9.850 2.810 ;
        RECT  9.545 2.605 9.785 2.765 ;
        RECT  9.285 2.605 9.545 2.865 ;
        RECT  9.505 0.695 9.510 0.870 ;
        RECT  9.245 0.610 9.505 0.870 ;
        END
        ANTENNADIFFAREA     0.2231 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.195 1.035 10.455 2.445 ;
        END
        ANTENNADIFFAREA     0.2156 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.265 1.735 1.525 ;
        RECT  1.690 1.265 1.715 2.400 ;
        RECT  1.505 1.265 1.690 2.430 ;
        RECT  1.475 1.265 1.505 1.525 ;
        RECT  1.475 2.270 1.505 2.430 ;
        RECT  1.215 2.270 1.475 2.530 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.740 4.250 2.035 ;
        RECT  3.805 1.700 4.015 2.035 ;
        RECT  3.765 1.740 3.805 2.035 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.015 -0.250 10.580 0.250 ;
        RECT  9.755 -0.250 10.015 0.405 ;
        RECT  8.935 -0.250 9.755 0.250 ;
        RECT  8.675 -0.250 8.935 0.795 ;
        RECT  5.235 -0.250 8.675 0.250 ;
        RECT  4.975 -0.250 5.235 0.405 ;
        RECT  4.035 -0.250 4.975 0.250 ;
        RECT  3.775 -0.250 4.035 0.405 ;
        RECT  1.540 -0.250 3.775 0.250 ;
        RECT  1.280 -0.250 1.540 0.405 ;
        RECT  0.265 -0.250 1.280 0.250 ;
        RECT  0.265 1.035 0.385 1.295 ;
        RECT  0.105 -0.250 0.265 1.295 ;
        RECT  0.000 -0.250 0.105 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.055 3.440 10.580 3.940 ;
        RECT  9.795 3.285 10.055 3.940 ;
        RECT  8.975 3.440 9.795 3.940 ;
        RECT  8.715 2.895 8.975 3.940 ;
        RECT  7.220 3.440 8.715 3.940 ;
        RECT  6.960 2.985 7.220 3.940 ;
        RECT  5.310 3.440 6.960 3.940 ;
        RECT  5.050 3.105 5.310 3.940 ;
        RECT  4.035 3.440 5.050 3.940 ;
        RECT  3.775 3.105 4.035 3.940 ;
        RECT  1.675 3.440 3.775 3.940 ;
        RECT  1.415 3.285 1.675 3.940 ;
        RECT  0.385 3.440 1.415 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.545 1.120 9.670 2.340 ;
        RECT  9.510 1.120 9.545 2.345 ;
        RECT  9.295 1.120 9.510 1.380 ;
        RECT  9.285 2.085 9.510 2.345 ;
        RECT  8.630 2.170 9.285 2.330 ;
        RECT  8.925 1.175 9.085 1.600 ;
        RECT  7.835 1.175 8.925 1.335 ;
        RECT  8.370 2.170 8.630 2.430 ;
        RECT  8.295 0.690 8.395 0.950 ;
        RECT  8.135 0.470 8.295 0.950 ;
        RECT  5.575 0.470 8.135 0.630 ;
        RECT  7.810 0.935 7.835 2.795 ;
        RECT  7.675 0.935 7.810 2.895 ;
        RECT  7.445 0.935 7.675 1.100 ;
        RECT  7.550 2.635 7.675 2.895 ;
        RECT  7.125 2.635 7.550 2.795 ;
        RECT  7.335 1.280 7.495 2.340 ;
        RECT  7.185 0.840 7.445 1.100 ;
        RECT  6.775 1.280 7.335 1.440 ;
        RECT  6.965 2.085 7.125 2.795 ;
        RECT  6.615 0.810 6.875 1.100 ;
        RECT  6.615 1.280 6.775 3.220 ;
        RECT  5.925 0.810 6.615 0.970 ;
        RECT  6.365 1.280 6.615 1.440 ;
        RECT  5.880 3.060 6.615 3.220 ;
        RECT  6.275 1.695 6.435 2.845 ;
        RECT  6.105 1.150 6.365 1.440 ;
        RECT  5.925 1.695 6.275 1.855 ;
        RECT  5.280 2.040 6.020 2.200 ;
        RECT  5.765 0.810 5.925 1.855 ;
        RECT  5.670 2.380 5.880 3.220 ;
        RECT  4.740 1.690 5.765 1.850 ;
        RECT  5.620 2.380 5.670 2.640 ;
        RECT  5.415 0.470 5.575 1.190 ;
        RECT  5.255 1.030 5.415 1.190 ;
        RECT  5.120 2.040 5.280 2.890 ;
        RECT  4.995 1.030 5.255 1.290 ;
        RECT  4.615 2.730 5.120 2.890 ;
        RECT  3.185 2.390 4.940 2.550 ;
        RECT  4.665 1.690 4.740 2.165 ;
        RECT  4.505 1.030 4.665 2.165 ;
        RECT  4.365 0.520 4.625 0.780 ;
        RECT  4.355 2.730 4.615 2.990 ;
        RECT  4.405 1.030 4.505 1.505 ;
        RECT  4.480 2.005 4.505 2.165 ;
        RECT  3.655 1.345 4.405 1.505 ;
        RECT  2.845 0.585 4.365 0.745 ;
        RECT  3.435 2.730 4.355 2.890 ;
        RECT  3.175 2.730 3.435 2.990 ;
        RECT  3.025 0.925 3.185 2.550 ;
        RECT  2.845 2.730 3.175 2.890 ;
        RECT  2.685 0.585 2.845 2.890 ;
        RECT  2.345 0.430 2.505 2.870 ;
        RECT  0.605 0.585 2.345 0.745 ;
        RECT  0.795 2.710 2.345 2.870 ;
        RECT  2.005 0.925 2.165 1.410 ;
        RECT  0.970 0.925 2.005 1.085 ;
        RECT  0.825 0.925 0.970 1.295 ;
        RECT  0.665 0.925 0.825 2.305 ;
        RECT  0.535 2.660 0.795 2.920 ;
        RECT  0.445 0.430 0.605 0.745 ;
    END
END SDFFSXL

MACRO SDFFRX4
    CLASS CORE ;
    FOREIGN SDFFRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.640 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.450 1.970 4.015 2.400 ;
        END
        ANTENNAGATEAREA     0.1456 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.350 1.955 2.450 2.215 ;
        RECT  2.190 1.955 2.350 2.340 ;
        RECT  0.880 2.180 2.190 2.340 ;
        RECT  0.795 2.180 0.880 2.480 ;
        RECT  0.585 2.110 0.795 2.480 ;
        RECT  0.570 2.220 0.585 2.480 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.650 1.480 12.290 1.640 ;
        RECT  11.580 1.290 11.650 1.640 ;
        RECT  11.420 0.470 11.580 1.640 ;
        RECT  8.430 0.470 11.420 0.630 ;
        RECT  8.420 0.470 8.430 0.695 ;
        RECT  8.260 0.470 8.420 1.040 ;
        RECT  8.155 0.880 8.260 1.040 ;
        RECT  8.130 0.880 8.155 1.170 ;
        RECT  7.790 0.880 8.130 1.430 ;
        RECT  7.720 0.880 7.790 1.040 ;
        RECT  7.560 0.470 7.720 1.040 ;
        RECT  5.655 0.470 7.560 0.630 ;
        RECT  5.495 0.470 5.655 0.745 ;
        RECT  4.345 0.585 5.495 0.745 ;
        RECT  4.185 0.585 4.345 1.380 ;
        RECT  4.015 1.220 4.185 1.380 ;
        RECT  3.755 1.220 4.015 1.545 ;
        END
        ANTENNAGATEAREA     0.4355 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.875 0.620 13.895 1.220 ;
        RECT  13.730 0.620 13.875 1.555 ;
        RECT  13.635 0.620 13.730 2.335 ;
        RECT  13.470 1.105 13.635 2.335 ;
        RECT  13.465 1.105 13.470 1.990 ;
        END
        ANTENNADIFFAREA     0.8312 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.655 0.675 14.915 1.275 ;
        RECT  14.625 1.975 14.840 2.335 ;
        RECT  14.625 1.035 14.655 1.275 ;
        RECT  14.580 1.035 14.625 2.335 ;
        RECT  14.385 1.035 14.580 2.215 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.665 1.535 1.925 ;
        RECT  1.045 1.665 1.255 1.990 ;
        RECT  0.955 1.665 1.045 1.925 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.575 4.745 1.925 ;
        RECT  4.380 1.575 4.475 1.990 ;
        RECT  4.265 1.700 4.380 1.990 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.425 -0.250 15.640 0.250 ;
        RECT  15.165 -0.250 15.425 1.265 ;
        RECT  14.405 -0.250 15.165 0.250 ;
        RECT  14.145 -0.250 14.405 0.775 ;
        RECT  13.350 -0.250 14.145 0.250 ;
        RECT  13.090 -0.250 13.350 0.405 ;
        RECT  12.040 -0.250 13.090 0.250 ;
        RECT  11.780 -0.250 12.040 0.405 ;
        RECT  8.060 -0.250 11.780 0.250 ;
        RECT  7.900 -0.250 8.060 0.625 ;
        RECT  5.310 -0.250 7.900 0.250 ;
        RECT  5.050 -0.250 5.310 0.405 ;
        RECT  3.545 -0.250 5.050 0.250 ;
        RECT  3.285 -0.250 3.545 0.690 ;
        RECT  0.385 -0.250 3.285 0.250 ;
        RECT  0.125 -0.250 0.385 0.845 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.390 3.440 15.640 3.940 ;
        RECT  15.130 2.895 15.390 3.940 ;
        RECT  14.270 3.405 15.130 3.940 ;
        RECT  14.010 2.895 14.270 3.940 ;
        RECT  13.160 3.405 14.010 3.940 ;
        RECT  12.900 2.895 13.160 3.940 ;
        RECT  11.990 3.405 12.900 3.940 ;
        RECT  11.730 3.285 11.990 3.940 ;
        RECT  9.205 3.405 11.730 3.940 ;
        RECT  8.945 2.975 9.205 3.940 ;
        RECT  7.870 3.440 8.945 3.940 ;
        RECT  7.710 2.560 7.870 3.940 ;
        RECT  7.335 3.440 7.710 3.940 ;
        RECT  7.075 2.800 7.335 3.940 ;
        RECT  4.955 3.440 7.075 3.940 ;
        RECT  4.695 3.285 4.955 3.940 ;
        RECT  3.735 3.440 4.695 3.940 ;
        RECT  3.475 2.945 3.735 3.940 ;
        RECT  1.350 3.440 3.475 3.940 ;
        RECT  1.090 2.600 1.350 3.940 ;
        RECT  0.000 3.440 1.090 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.115 1.560 15.185 2.675 ;
        RECT  15.025 1.510 15.115 2.675 ;
        RECT  14.855 1.510 15.025 1.770 ;
        RECT  13.155 2.515 15.025 2.675 ;
        RECT  12.995 0.915 13.155 2.675 ;
        RECT  12.940 0.915 12.995 1.995 ;
        RECT  12.580 2.515 12.995 2.675 ;
        RECT  12.925 0.695 12.940 1.995 ;
        RECT  12.680 0.695 12.925 1.295 ;
        RECT  11.450 1.835 12.925 1.995 ;
        RECT  11.240 2.175 12.815 2.335 ;
        RECT  12.320 2.515 12.580 3.195 ;
        RECT  11.155 2.965 11.415 3.225 ;
        RECT  11.080 0.810 11.240 2.785 ;
        RECT  9.635 2.965 11.155 3.125 ;
        RECT  10.240 0.810 11.080 0.970 ;
        RECT  10.950 2.525 11.080 2.785 ;
        RECT  10.190 2.625 10.950 2.785 ;
        RECT  10.650 1.150 10.780 1.310 ;
        RECT  10.650 2.255 10.700 2.415 ;
        RECT  10.490 1.150 10.650 2.415 ;
        RECT  8.770 1.650 10.490 1.810 ;
        RECT  10.440 2.255 10.490 2.415 ;
        RECT  9.980 0.810 10.240 1.070 ;
        RECT  9.930 2.500 10.190 2.785 ;
        RECT  9.630 0.810 9.730 1.070 ;
        RECT  8.555 2.285 9.680 2.445 ;
        RECT  9.475 2.625 9.635 3.125 ;
        RECT  9.470 0.810 9.630 1.295 ;
        RECT  8.210 2.625 9.475 2.785 ;
        RECT  8.770 1.135 9.470 1.295 ;
        RECT  8.610 1.135 8.770 1.810 ;
        RECT  8.555 1.650 8.610 1.810 ;
        RECT  8.395 1.650 8.555 2.445 ;
        RECT  7.820 1.650 8.395 1.810 ;
        RECT  8.050 2.090 8.210 2.785 ;
        RECT  7.380 2.090 8.050 2.250 ;
        RECT  7.560 1.650 7.820 1.910 ;
        RECT  6.835 2.430 7.495 2.590 ;
        RECT  7.220 0.810 7.380 2.250 ;
        RECT  6.015 0.810 7.220 0.970 ;
        RECT  6.835 1.150 7.035 1.310 ;
        RECT  6.675 1.150 6.835 2.930 ;
        RECT  6.335 2.770 6.675 2.930 ;
        RECT  6.415 1.150 6.465 1.310 ;
        RECT  6.255 1.150 6.415 2.555 ;
        RECT  6.175 2.770 6.335 3.105 ;
        RECT  6.205 1.150 6.255 1.310 ;
        RECT  5.875 2.395 6.255 2.555 ;
        RECT  4.135 2.945 6.175 3.105 ;
        RECT  6.015 1.555 6.075 1.815 ;
        RECT  5.975 0.810 6.015 1.815 ;
        RECT  5.855 0.810 5.975 2.160 ;
        RECT  5.715 2.395 5.875 2.765 ;
        RECT  5.630 0.970 5.855 1.230 ;
        RECT  5.815 1.555 5.855 2.160 ;
        RECT  5.455 2.000 5.815 2.160 ;
        RECT  3.270 2.605 5.715 2.765 ;
        RECT  5.515 1.450 5.565 1.710 ;
        RECT  5.310 1.450 5.515 1.815 ;
        RECT  5.295 2.000 5.455 2.295 ;
        RECT  5.150 1.030 5.310 1.815 ;
        RECT  4.790 1.030 5.150 1.190 ;
        RECT  5.110 1.655 5.150 1.815 ;
        RECT  4.950 1.655 5.110 2.375 ;
        RECT  4.210 2.215 4.950 2.375 ;
        RECT  4.530 0.930 4.790 1.190 ;
        RECT  3.845 0.560 4.005 1.035 ;
        RECT  3.035 0.875 3.845 1.035 ;
        RECT  3.110 1.215 3.270 2.765 ;
        RECT  2.355 1.215 3.110 1.375 ;
        RECT  2.625 2.605 3.110 2.765 ;
        RECT  2.935 0.775 3.035 1.035 ;
        RECT  2.775 0.480 2.935 1.035 ;
        RECT  2.830 1.955 2.930 2.215 ;
        RECT  2.670 1.565 2.830 2.215 ;
        RECT  1.360 0.480 2.775 0.640 ;
        RECT  2.015 1.565 2.670 1.725 ;
        RECT  2.025 2.535 2.625 2.795 ;
        RECT  2.195 0.855 2.355 1.375 ;
        RECT  1.925 0.855 2.195 1.015 ;
        RECT  1.855 1.265 2.015 1.725 ;
        RECT  1.755 1.265 1.855 1.605 ;
        RECT  0.965 1.265 1.755 1.425 ;
        RECT  1.100 0.480 1.360 0.755 ;
        RECT  0.705 1.030 0.965 1.425 ;
        RECT  0.365 1.265 0.705 1.425 ;
        RECT  0.420 2.720 0.680 2.980 ;
        RECT  0.365 2.720 0.420 2.880 ;
        RECT  0.205 1.265 0.365 2.880 ;
    END
END SDFFRX4

MACRO SDFFRX2
    CLASS CORE ;
    FOREIGN SDFFRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.420 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.820 1.955 3.100 2.400 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.560 1.645 1.820 1.905 ;
        RECT  1.255 1.745 1.560 1.905 ;
        RECT  1.045 1.700 1.255 1.990 ;
        RECT  0.885 1.700 1.045 1.940 ;
        RECT  0.625 1.680 0.885 1.940 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.295 1.405 9.555 1.665 ;
        RECT  8.910 1.405 9.295 1.565 ;
        RECT  8.750 0.470 8.910 1.565 ;
        RECT  7.635 0.470 8.750 0.630 ;
        RECT  7.475 0.470 7.635 1.330 ;
        RECT  7.285 1.170 7.475 1.330 ;
        RECT  7.025 1.170 7.285 1.430 ;
        RECT  6.955 1.170 7.025 1.330 ;
        RECT  6.795 0.470 6.955 1.330 ;
        RECT  4.890 0.470 6.795 0.630 ;
        RECT  4.730 0.470 4.890 0.745 ;
        RECT  3.545 0.585 4.730 0.745 ;
        RECT  3.545 1.700 3.555 1.990 ;
        RECT  3.385 0.585 3.545 1.990 ;
        RECT  3.345 1.400 3.385 1.990 ;
        RECT  3.115 1.400 3.345 1.660 ;
        END
        ANTENNAGATEAREA     0.2444 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.840 1.105 10.915 2.755 ;
        RECT  10.630 0.515 10.840 2.755 ;
        RECT  10.480 0.515 10.630 0.775 ;
        END
        ANTENNADIFFAREA     0.5026 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.650 2.155 11.865 2.755 ;
        RECT  11.465 0.845 11.760 1.105 ;
        RECT  11.605 2.110 11.650 2.755 ;
        RECT  11.465 2.110 11.605 2.315 ;
        RECT  11.350 0.845 11.465 2.315 ;
        RECT  11.305 0.945 11.350 2.315 ;
        RECT  11.165 1.105 11.305 1.765 ;
        END
        ANTENNADIFFAREA     0.4028 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.930 1.715 3.220 ;
        RECT  1.340 2.930 1.505 3.180 ;
        RECT  1.080 2.920 1.340 3.180 ;
        END
        ANTENNAGATEAREA     0.1443 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.050 1.495 4.310 1.755 ;
        RECT  4.015 1.495 4.050 1.655 ;
        RECT  3.805 1.290 4.015 1.655 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.270 -0.250 12.420 0.250 ;
        RECT  12.010 -0.250 12.270 1.095 ;
        RECT  11.310 -0.250 12.010 0.250 ;
        RECT  11.050 -0.250 11.310 0.405 ;
        RECT  9.455 -0.250 11.050 0.250 ;
        RECT  9.195 -0.250 9.455 1.135 ;
        RECT  7.295 -0.250 9.195 0.250 ;
        RECT  7.135 -0.250 7.295 0.625 ;
        RECT  4.545 -0.250 7.135 0.250 ;
        RECT  4.285 -0.250 4.545 0.405 ;
        RECT  3.755 -0.250 4.285 0.250 ;
        RECT  3.495 -0.250 3.755 0.405 ;
        RECT  0.455 -0.250 3.495 0.250 ;
        RECT  0.195 -0.250 0.455 0.845 ;
        RECT  0.000 -0.250 0.195 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.265 3.440 12.420 3.940 ;
        RECT  12.005 3.285 12.265 3.940 ;
        RECT  11.290 3.440 12.005 3.940 ;
        RECT  10.690 3.285 11.290 3.940 ;
        RECT  9.120 3.440 10.690 3.940 ;
        RECT  8.860 3.285 9.120 3.940 ;
        RECT  7.085 3.440 8.860 3.940 ;
        RECT  6.925 2.560 7.085 3.940 ;
        RECT  6.560 3.440 6.925 3.940 ;
        RECT  6.300 2.800 6.560 3.940 ;
        RECT  4.530 3.440 6.300 3.940 ;
        RECT  4.270 3.285 4.530 3.940 ;
        RECT  3.105 3.440 4.270 3.940 ;
        RECT  2.845 2.945 3.105 3.940 ;
        RECT  0.850 3.440 2.845 3.940 ;
        RECT  0.900 2.335 1.160 2.595 ;
        RECT  0.850 2.435 0.900 2.595 ;
        RECT  0.690 2.435 0.850 3.940 ;
        RECT  0.000 3.440 0.690 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.065 1.725 12.225 3.105 ;
        RECT  12.010 1.725 12.065 1.885 ;
        RECT  10.330 2.945 12.065 3.105 ;
        RECT  11.750 1.625 12.010 1.885 ;
        RECT  10.320 1.035 10.330 3.105 ;
        RECT  10.160 1.035 10.320 3.110 ;
        RECT  10.045 1.035 10.160 2.010 ;
        RECT  9.745 2.950 10.160 3.110 ;
        RECT  9.055 1.850 10.045 2.010 ;
        RECT  9.720 2.285 9.980 2.565 ;
        RECT  9.485 2.950 9.745 3.210 ;
        RECT  8.465 2.285 9.720 2.445 ;
        RECT  8.795 1.750 9.055 2.010 ;
        RECT  8.320 2.980 8.580 3.240 ;
        RECT  8.465 0.810 8.565 1.070 ;
        RECT  8.305 0.810 8.465 2.665 ;
        RECT  7.425 3.015 8.320 3.175 ;
        RECT  8.115 2.065 8.305 2.665 ;
        RECT  7.865 0.820 8.005 1.860 ;
        RECT  7.845 0.820 7.865 2.835 ;
        RECT  7.605 1.700 7.845 2.835 ;
        RECT  6.960 1.700 7.605 1.860 ;
        RECT  7.265 2.090 7.425 3.175 ;
        RECT  6.615 2.090 7.265 2.250 ;
        RECT  6.800 1.650 6.960 1.910 ;
        RECT  6.070 2.430 6.730 2.590 ;
        RECT  6.455 0.810 6.615 2.250 ;
        RECT  5.230 0.810 6.455 0.970 ;
        RECT  6.070 1.150 6.270 1.310 ;
        RECT  5.910 1.150 6.070 2.930 ;
        RECT  5.580 2.770 5.910 2.930 ;
        RECT  5.650 1.150 5.700 1.310 ;
        RECT  5.490 1.150 5.650 2.585 ;
        RECT  5.420 2.770 5.580 3.105 ;
        RECT  5.440 1.150 5.490 1.310 ;
        RECT  5.110 2.425 5.490 2.585 ;
        RECT  3.505 2.945 5.420 3.105 ;
        RECT  5.230 1.555 5.290 1.815 ;
        RECT  5.190 0.810 5.230 1.815 ;
        RECT  5.070 0.810 5.190 2.235 ;
        RECT  4.950 2.425 5.110 2.765 ;
        RECT  4.865 0.945 5.070 1.205 ;
        RECT  5.030 1.555 5.070 2.235 ;
        RECT  4.850 2.075 5.030 2.235 ;
        RECT  2.610 2.605 4.950 2.765 ;
        RECT  4.660 1.450 4.800 1.710 ;
        RECT  4.500 0.945 4.660 2.175 ;
        RECT  3.855 0.945 4.500 1.105 ;
        RECT  4.100 2.015 4.500 2.175 ;
        RECT  3.840 2.015 4.100 2.275 ;
        RECT  3.155 0.600 3.205 1.200 ;
        RECT  2.945 0.480 3.155 1.200 ;
        RECT  1.415 0.480 2.945 0.640 ;
        RECT  2.450 0.830 2.610 2.765 ;
        RECT  2.035 0.830 2.450 0.990 ;
        RECT  2.030 2.395 2.450 2.555 ;
        RECT  2.090 1.210 2.250 2.215 ;
        RECT  1.035 1.210 2.090 1.370 ;
        RECT  1.770 2.395 2.030 2.655 ;
        RECT  1.155 0.480 1.415 0.755 ;
        RECT  0.775 1.030 1.035 1.370 ;
        RECT  0.410 1.210 0.775 1.370 ;
        RECT  0.410 2.180 0.510 2.440 ;
        RECT  0.250 1.210 0.410 2.440 ;
    END
END SDFFRX2

MACRO SDFFRX1
    CLASS CORE ;
    FOREIGN SDFFRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 2.930 2.305 3.240 ;
        RECT  1.965 2.930 2.045 3.220 ;
        RECT  1.805 2.930 1.965 3.180 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.750 1.585 2.010 ;
        RECT  0.795 1.750 1.230 1.910 ;
        RECT  0.755 1.700 0.795 1.990 ;
        RECT  0.585 1.680 0.755 1.990 ;
        RECT  0.495 1.680 0.585 1.940 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.445 9.105 1.745 ;
        RECT  8.840 1.445 9.100 1.795 ;
        RECT  8.450 1.445 8.840 1.605 ;
        RECT  8.290 0.470 8.450 1.605 ;
        RECT  7.170 0.470 8.290 0.630 ;
        RECT  7.010 0.470 7.170 1.330 ;
        RECT  6.825 1.170 7.010 1.330 ;
        RECT  6.565 1.170 6.825 1.430 ;
        RECT  6.490 1.170 6.565 1.330 ;
        RECT  6.330 0.470 6.490 1.330 ;
        RECT  4.430 0.470 6.330 0.630 ;
        RECT  4.270 0.470 4.430 0.745 ;
        RECT  3.095 0.585 4.270 0.745 ;
        RECT  2.910 0.585 3.095 1.990 ;
        RECT  2.885 1.105 2.910 1.990 ;
        RECT  2.655 1.400 2.885 1.660 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.260 1.700 10.455 1.990 ;
        RECT  10.100 0.690 10.260 2.315 ;
        RECT  9.890 0.690 10.100 0.850 ;
        RECT  9.970 2.110 10.100 2.315 ;
        RECT  9.940 2.155 9.970 2.315 ;
        RECT  9.680 2.155 9.940 2.755 ;
        RECT  9.630 0.590 9.890 0.850 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.910 1.105 10.915 2.755 ;
        RECT  10.705 0.845 10.910 2.755 ;
        RECT  10.650 0.845 10.705 1.105 ;
        RECT  10.655 2.155 10.705 2.755 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 2.535 1.275 3.180 ;
        RECT  1.045 2.520 1.255 3.180 ;
        RECT  1.015 2.535 1.045 3.180 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.495 3.850 1.755 ;
        RECT  3.555 1.495 3.590 1.655 ;
        RECT  3.345 1.290 3.555 1.655 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.460 -0.250 11.040 0.250 ;
        RECT  10.200 -0.250 10.460 0.405 ;
        RECT  8.980 -0.250 10.200 0.250 ;
        RECT  8.720 -0.250 8.980 1.145 ;
        RECT  6.830 -0.250 8.720 0.250 ;
        RECT  6.670 -0.250 6.830 0.625 ;
        RECT  4.085 -0.250 6.670 0.250 ;
        RECT  3.825 -0.250 4.085 0.405 ;
        RECT  3.145 -0.250 3.825 0.250 ;
        RECT  2.885 -0.250 3.145 0.405 ;
        RECT  0.385 -0.250 2.885 0.250 ;
        RECT  0.125 -0.250 0.385 1.055 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.340 3.440 11.040 3.940 ;
        RECT  9.740 3.285 10.340 3.940 ;
        RECT  8.300 3.440 9.740 3.940 ;
        RECT  8.040 3.285 8.300 3.940 ;
        RECT  6.110 3.440 8.040 3.940 ;
        RECT  5.850 2.800 6.110 3.940 ;
        RECT  4.070 3.440 5.850 3.940 ;
        RECT  3.810 3.285 4.070 3.940 ;
        RECT  2.755 3.440 3.810 3.940 ;
        RECT  2.495 2.895 2.755 3.940 ;
        RECT  0.820 3.440 2.495 3.940 ;
        RECT  0.560 2.895 0.820 3.940 ;
        RECT  0.000 3.440 0.560 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.500 2.945 10.730 3.105 ;
        RECT  9.600 1.130 9.860 1.390 ;
        RECT  9.500 1.180 9.600 1.390 ;
        RECT  9.340 1.180 9.500 3.160 ;
        RECT  8.510 1.980 9.340 2.140 ;
        RECT  8.665 3.000 9.340 3.160 ;
        RECT  8.900 2.550 9.160 2.790 ;
        RECT  8.050 2.550 8.900 2.710 ;
        RECT  8.250 1.785 8.510 2.140 ;
        RECT  8.050 0.820 8.100 0.980 ;
        RECT  7.890 0.820 8.050 2.710 ;
        RECT  7.840 0.820 7.890 0.980 ;
        RECT  7.555 2.500 7.890 2.710 ;
        RECT  7.500 2.980 7.760 3.240 ;
        RECT  7.295 2.500 7.555 2.760 ;
        RECT  7.350 0.820 7.510 1.910 ;
        RECT  6.605 2.980 7.500 3.140 ;
        RECT  6.995 1.750 7.350 1.910 ;
        RECT  6.995 2.510 7.045 2.770 ;
        RECT  6.835 1.750 6.995 2.770 ;
        RECT  6.590 1.750 6.835 1.910 ;
        RECT  6.785 2.510 6.835 2.770 ;
        RECT  6.445 2.090 6.605 3.140 ;
        RECT  6.330 1.650 6.590 1.910 ;
        RECT  6.150 2.090 6.445 2.250 ;
        RECT  5.610 2.430 6.265 2.590 ;
        RECT  5.990 0.810 6.150 2.250 ;
        RECT  4.790 0.810 5.990 0.970 ;
        RECT  5.610 1.150 5.810 1.310 ;
        RECT  5.450 1.150 5.610 2.930 ;
        RECT  5.215 2.770 5.450 2.930 ;
        RECT  5.190 1.150 5.240 1.310 ;
        RECT  4.960 2.770 5.215 3.105 ;
        RECT  5.030 1.150 5.190 2.585 ;
        RECT  4.980 1.150 5.030 1.310 ;
        RECT  4.650 2.425 5.030 2.585 ;
        RECT  3.265 2.945 4.960 3.105 ;
        RECT  4.790 1.555 4.820 1.815 ;
        RECT  4.720 0.810 4.790 1.815 ;
        RECT  4.650 0.810 4.720 2.170 ;
        RECT  4.630 0.810 4.650 2.235 ;
        RECT  4.390 2.425 4.650 2.765 ;
        RECT  4.405 0.945 4.630 1.205 ;
        RECT  4.560 1.555 4.630 2.235 ;
        RECT  4.390 2.010 4.560 2.235 ;
        RECT  3.610 2.605 4.390 2.765 ;
        RECT  4.200 1.450 4.340 1.710 ;
        RECT  4.040 0.945 4.200 2.130 ;
        RECT  3.395 0.945 4.040 1.105 ;
        RECT  3.640 1.970 4.040 2.130 ;
        RECT  3.380 1.970 3.640 2.230 ;
        RECT  3.450 2.435 3.610 2.765 ;
        RECT  2.355 2.435 3.450 2.595 ;
        RECT  2.995 2.800 3.265 3.105 ;
        RECT  2.535 0.515 2.695 1.220 ;
        RECT  0.955 0.515 2.535 0.675 ;
        RECT  2.350 1.640 2.355 2.595 ;
        RECT  2.195 0.910 2.350 2.595 ;
        RECT  2.190 0.910 2.195 1.800 ;
        RECT  1.535 2.435 2.195 2.595 ;
        RECT  1.835 0.910 2.190 1.070 ;
        RECT  1.990 1.990 2.015 2.250 ;
        RECT  1.830 1.250 1.990 2.250 ;
        RECT  1.575 0.860 1.835 1.070 ;
        RECT  0.955 1.250 1.830 1.410 ;
        RECT  0.695 0.515 0.955 0.785 ;
        RECT  0.695 1.035 0.955 1.410 ;
        RECT  0.285 1.250 0.695 1.410 ;
        RECT  0.285 2.180 0.385 2.440 ;
        RECT  0.125 1.250 0.285 2.440 ;
    END
END SDFFRX1

MACRO SDFFRXL
    CLASS CORE ;
    FOREIGN SDFFRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 2.930 2.305 3.240 ;
        RECT  1.965 2.930 2.045 3.220 ;
        RECT  1.805 2.930 1.965 3.180 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.750 1.585 2.010 ;
        RECT  0.795 1.780 1.230 1.940 ;
        RECT  0.755 1.700 0.795 1.990 ;
        RECT  0.585 1.680 0.755 1.990 ;
        RECT  0.495 1.680 0.585 1.940 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.900 1.480 9.160 1.795 ;
        RECT  8.615 1.480 8.900 1.640 ;
        RECT  8.495 1.105 8.615 1.640 ;
        RECT  8.335 0.470 8.495 1.640 ;
        RECT  7.175 0.470 8.335 0.630 ;
        RECT  7.015 0.470 7.175 1.330 ;
        RECT  6.825 1.170 7.015 1.330 ;
        RECT  6.565 1.170 6.825 1.430 ;
        RECT  6.495 1.170 6.565 1.330 ;
        RECT  6.335 0.470 6.495 1.330 ;
        RECT  4.430 0.470 6.335 0.630 ;
        RECT  4.270 0.470 4.430 0.745 ;
        RECT  3.095 0.585 4.270 0.745 ;
        RECT  2.910 0.585 3.095 1.990 ;
        RECT  2.885 1.105 2.910 1.990 ;
        RECT  2.655 1.400 2.885 1.660 ;
        END
        ANTENNAGATEAREA     0.1274 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.260 1.700 10.455 1.990 ;
        RECT  10.100 0.695 10.260 2.315 ;
        RECT  9.860 0.695 10.100 0.855 ;
        RECT  9.970 2.110 10.100 2.315 ;
        RECT  9.890 2.155 9.970 2.315 ;
        RECT  9.730 2.155 9.890 2.585 ;
        RECT  9.600 0.595 9.860 0.855 ;
        END
        ANTENNADIFFAREA     0.2142 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.910 1.105 10.915 2.585 ;
        RECT  10.705 0.845 10.910 2.585 ;
        RECT  10.650 0.845 10.705 1.105 ;
        RECT  10.655 2.325 10.705 2.585 ;
        END
        ANTENNADIFFAREA     0.2142 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 2.535 1.275 3.180 ;
        RECT  1.045 2.520 1.255 3.180 ;
        RECT  1.015 2.535 1.045 3.180 ;
        END
        ANTENNAGATEAREA     0.0650 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.495 3.850 1.755 ;
        RECT  3.555 1.495 3.590 1.655 ;
        RECT  3.345 1.290 3.555 1.655 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.460 -0.250 11.040 0.250 ;
        RECT  10.200 -0.250 10.460 0.405 ;
        RECT  9.035 -0.250 10.200 0.250 ;
        RECT  8.775 -0.250 9.035 0.800 ;
        RECT  6.835 -0.250 8.775 0.250 ;
        RECT  6.675 -0.250 6.835 0.625 ;
        RECT  4.085 -0.250 6.675 0.250 ;
        RECT  3.825 -0.250 4.085 0.405 ;
        RECT  3.145 -0.250 3.825 0.250 ;
        RECT  2.885 -0.250 3.145 0.405 ;
        RECT  0.385 -0.250 2.885 0.250 ;
        RECT  0.125 -0.250 0.385 1.055 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.340 3.440 11.040 3.940 ;
        RECT  9.740 3.285 10.340 3.940 ;
        RECT  8.355 3.440 9.740 3.940 ;
        RECT  8.095 3.285 8.355 3.940 ;
        RECT  6.110 3.440 8.095 3.940 ;
        RECT  5.850 2.775 6.110 3.940 ;
        RECT  4.070 3.440 5.850 3.940 ;
        RECT  3.810 3.285 4.070 3.940 ;
        RECT  2.755 3.440 3.810 3.940 ;
        RECT  2.495 2.895 2.755 3.940 ;
        RECT  0.820 3.440 2.495 3.940 ;
        RECT  0.560 2.895 0.820 3.940 ;
        RECT  0.000 3.440 0.560 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.545 2.945 10.745 3.105 ;
        RECT  9.545 1.130 9.845 1.390 ;
        RECT  9.540 1.130 9.545 3.105 ;
        RECT  9.380 1.130 9.540 3.160 ;
        RECT  8.580 1.975 9.380 2.135 ;
        RECT  8.685 3.000 9.380 3.160 ;
        RECT  8.935 2.550 9.195 2.790 ;
        RECT  8.045 2.550 8.935 2.710 ;
        RECT  8.315 1.835 8.580 2.135 ;
        RECT  8.045 0.825 8.145 1.085 ;
        RECT  7.885 0.825 8.045 2.710 ;
        RECT  7.590 2.500 7.885 2.710 ;
        RECT  7.530 2.980 7.790 3.240 ;
        RECT  7.330 2.500 7.590 2.760 ;
        RECT  6.580 2.980 7.530 3.140 ;
        RECT  7.360 0.825 7.520 1.860 ;
        RECT  7.020 1.700 7.360 1.860 ;
        RECT  6.860 1.700 7.020 2.775 ;
        RECT  6.590 1.700 6.860 1.860 ;
        RECT  6.760 2.515 6.860 2.775 ;
        RECT  6.330 1.650 6.590 1.910 ;
        RECT  6.420 2.090 6.580 3.140 ;
        RECT  6.150 2.090 6.420 2.250 ;
        RECT  5.610 2.430 6.210 2.590 ;
        RECT  5.990 0.810 6.150 2.250 ;
        RECT  4.790 0.810 5.990 0.970 ;
        RECT  5.610 1.150 5.810 1.410 ;
        RECT  5.550 1.150 5.610 2.930 ;
        RECT  5.450 1.200 5.550 2.930 ;
        RECT  5.120 2.770 5.450 2.930 ;
        RECT  5.190 1.150 5.240 1.310 ;
        RECT  5.030 1.150 5.190 2.585 ;
        RECT  4.960 2.770 5.120 3.105 ;
        RECT  4.980 1.150 5.030 1.310 ;
        RECT  4.650 2.425 5.030 2.585 ;
        RECT  3.265 2.945 4.960 3.105 ;
        RECT  4.790 1.555 4.820 1.815 ;
        RECT  4.720 0.810 4.790 1.815 ;
        RECT  4.630 0.810 4.720 2.235 ;
        RECT  4.490 2.425 4.650 2.765 ;
        RECT  4.405 0.945 4.630 1.205 ;
        RECT  4.560 1.555 4.630 2.235 ;
        RECT  4.390 2.075 4.560 2.235 ;
        RECT  3.610 2.605 4.490 2.765 ;
        RECT  4.200 1.450 4.340 1.710 ;
        RECT  4.190 0.945 4.200 1.710 ;
        RECT  4.040 0.945 4.190 2.180 ;
        RECT  3.395 0.945 4.040 1.105 ;
        RECT  4.030 1.500 4.040 2.180 ;
        RECT  3.640 2.020 4.030 2.180 ;
        RECT  3.380 1.970 3.640 2.230 ;
        RECT  3.450 2.435 3.610 2.765 ;
        RECT  2.355 2.435 3.450 2.595 ;
        RECT  2.995 2.800 3.265 3.105 ;
        RECT  2.535 0.515 2.695 1.200 ;
        RECT  0.955 0.515 2.535 0.675 ;
        RECT  2.350 1.640 2.355 2.595 ;
        RECT  2.195 0.910 2.350 2.595 ;
        RECT  2.190 0.910 2.195 1.800 ;
        RECT  1.535 2.435 2.195 2.595 ;
        RECT  1.835 0.910 2.190 1.070 ;
        RECT  1.990 1.990 2.015 2.250 ;
        RECT  1.830 1.250 1.990 2.250 ;
        RECT  1.575 0.860 1.835 1.070 ;
        RECT  0.955 1.250 1.830 1.410 ;
        RECT  0.695 0.515 0.955 0.785 ;
        RECT  0.695 1.035 0.955 1.410 ;
        RECT  0.285 1.250 0.695 1.410 ;
        RECT  0.285 2.180 0.385 2.440 ;
        RECT  0.125 1.250 0.285 2.440 ;
    END
END SDFFRXL

MACRO SDFFQXL
    CLASS CORE ;
    FOREIGN SDFFQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.490 1.310 2.005 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.060 1.980 2.320 ;
        RECT  1.660 2.060 1.715 2.765 ;
        RECT  1.505 2.110 1.660 2.765 ;
        RECT  0.375 2.605 1.505 2.765 ;
        RECT  0.215 1.475 0.375 2.765 ;
        RECT  0.125 1.475 0.215 2.175 ;
        RECT  0.115 1.475 0.125 1.765 ;
        END
        ANTENNAGATEAREA     0.1196 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.600 2.745 8.615 3.025 ;
        RECT  8.440 0.520 8.600 3.025 ;
        RECT  8.155 0.520 8.440 0.780 ;
        RECT  8.405 2.745 8.440 3.025 ;
        RECT  7.970 2.765 8.405 3.025 ;
        RECT  7.970 0.470 8.155 0.780 ;
        RECT  7.945 0.470 7.970 0.760 ;
        RECT  7.920 0.500 7.945 0.760 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 1.290 2.175 1.580 ;
        RECT  1.965 1.290 2.145 1.840 ;
        RECT  1.840 1.580 1.965 1.840 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 2.110 4.595 2.400 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.655 -0.250 8.740 0.250 ;
        RECT  7.395 -0.250 7.655 0.405 ;
        RECT  6.035 -0.250 7.395 0.250 ;
        RECT  5.775 -0.250 6.035 1.005 ;
        RECT  4.440 -0.250 5.775 0.250 ;
        RECT  3.840 -0.250 4.440 0.625 ;
        RECT  1.690 -0.250 3.840 0.250 ;
        RECT  1.430 -0.250 1.690 0.405 ;
        RECT  0.360 -0.250 1.430 0.250 ;
        RECT  0.360 1.035 0.385 1.295 ;
        RECT  0.125 -0.250 0.360 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.685 3.440 8.740 3.940 ;
        RECT  7.425 2.555 7.685 3.940 ;
        RECT  5.860 3.440 7.425 3.940 ;
        RECT  5.600 3.285 5.860 3.940 ;
        RECT  4.850 3.440 5.600 3.940 ;
        RECT  4.590 3.285 4.850 3.940 ;
        RECT  3.950 3.440 4.590 3.940 ;
        RECT  3.690 3.285 3.950 3.940 ;
        RECT  1.865 3.440 3.690 3.940 ;
        RECT  1.605 3.285 1.865 3.940 ;
        RECT  0.385 3.440 1.605 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.100 1.035 8.260 2.320 ;
        RECT  7.975 1.035 8.100 1.295 ;
        RECT  8.000 2.055 8.100 2.320 ;
        RECT  7.400 2.055 8.000 2.215 ;
        RECT  7.740 1.495 7.905 1.755 ;
        RECT  7.580 1.240 7.740 1.755 ;
        RECT  6.940 1.240 7.580 1.400 ;
        RECT  7.240 1.590 7.400 2.215 ;
        RECT  7.140 1.590 7.240 1.850 ;
        RECT  6.855 0.455 7.115 0.715 ;
        RECT  6.935 0.935 6.940 1.400 ;
        RECT  6.775 0.935 6.935 2.690 ;
        RECT  6.405 0.555 6.855 0.715 ;
        RECT  6.630 0.935 6.775 1.095 ;
        RECT  6.720 2.530 6.775 2.690 ;
        RECT  6.460 2.530 6.720 2.790 ;
        RECT  6.455 2.040 6.595 2.300 ;
        RECT  6.405 1.305 6.455 2.300 ;
        RECT  6.295 0.555 6.405 2.300 ;
        RECT  6.245 0.555 6.295 1.465 ;
        RECT  6.190 2.140 6.295 2.300 ;
        RECT  5.845 1.305 6.245 1.465 ;
        RECT  6.030 2.140 6.190 3.105 ;
        RECT  5.855 1.685 6.115 1.945 ;
        RECT  4.420 2.945 6.030 3.105 ;
        RECT  5.845 1.785 5.855 1.945 ;
        RECT  5.685 1.205 5.845 1.465 ;
        RECT  5.685 1.785 5.845 2.750 ;
        RECT  4.980 2.590 5.685 2.750 ;
        RECT  5.345 0.595 5.505 2.290 ;
        RECT  5.120 0.595 5.345 0.855 ;
        RECT  5.170 2.030 5.345 2.290 ;
        RECT  5.005 1.105 5.165 1.365 ;
        RECT  5.005 0.595 5.120 0.755 ;
        RECT  4.845 0.430 5.005 0.755 ;
        RECT  4.980 1.205 5.005 1.365 ;
        RECT  4.820 1.205 4.980 2.750 ;
        RECT  4.745 0.430 4.845 0.590 ;
        RECT  3.630 1.715 4.820 1.875 ;
        RECT  2.900 1.375 4.420 1.535 ;
        RECT  4.160 2.580 4.420 3.105 ;
        RECT  4.015 0.935 4.275 1.195 ;
        RECT  3.165 2.940 4.160 3.105 ;
        RECT  3.490 0.935 4.015 1.095 ;
        RECT  3.370 1.715 3.630 1.975 ;
        RECT  3.330 0.770 3.490 1.095 ;
        RECT  2.560 0.770 3.330 0.930 ;
        RECT  3.060 2.710 3.165 3.105 ;
        RECT  2.900 2.370 3.070 2.530 ;
        RECT  3.005 2.710 3.060 3.100 ;
        RECT  2.560 2.710 3.005 2.870 ;
        RECT  2.740 1.110 2.900 2.530 ;
        RECT  2.220 3.050 2.670 3.210 ;
        RECT  2.400 0.770 2.560 2.870 ;
        RECT  2.220 0.430 2.480 0.590 ;
        RECT  2.370 1.270 2.400 1.530 ;
        RECT  2.060 0.430 2.220 0.775 ;
        RECT  2.060 2.945 2.220 3.210 ;
        RECT  0.800 0.615 2.060 0.775 ;
        RECT  0.965 2.945 2.060 3.105 ;
        RECT  1.580 1.090 1.740 1.350 ;
        RECT  0.955 1.090 1.580 1.250 ;
        RECT  0.855 2.265 1.185 2.425 ;
        RECT  0.705 2.945 0.965 3.205 ;
        RECT  0.855 1.035 0.955 1.295 ;
        RECT  0.695 1.035 0.855 2.425 ;
        RECT  0.540 0.455 0.800 0.775 ;
        RECT  0.555 1.955 0.695 2.215 ;
    END
END SDFFQXL

MACRO SDFFQX4
    CLASS CORE ;
    FOREIGN SDFFQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.490 1.310 2.005 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.220 1.980 2.380 ;
        RECT  1.505 2.110 1.715 2.685 ;
        RECT  0.375 2.525 1.505 2.685 ;
        RECT  0.215 1.475 0.375 2.685 ;
        RECT  0.125 1.475 0.215 2.175 ;
        RECT  0.115 1.475 0.125 1.765 ;
        END
        ANTENNAGATEAREA     0.1248 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.245 1.290 10.455 1.990 ;
        RECT  10.240 1.290 10.245 3.015 ;
        RECT  9.985 0.560 10.240 3.015 ;
        RECT  9.980 0.560 9.985 1.160 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 1.595 2.175 1.990 ;
        RECT  1.875 1.625 1.935 1.990 ;
        RECT  1.840 1.660 1.875 1.920 ;
        END
        ANTENNAGATEAREA     0.0897 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 2.110 4.310 2.400 ;
        END
        ANTENNAGATEAREA     0.1677 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.750 -0.250 11.040 0.250 ;
        RECT  10.490 -0.250 10.750 1.095 ;
        RECT  9.605 -0.250 10.490 0.250 ;
        RECT  9.345 -0.250 9.605 0.405 ;
        RECT  8.010 -0.250 9.345 0.250 ;
        RECT  7.750 -0.250 8.010 0.405 ;
        RECT  6.300 -0.250 7.750 0.250 ;
        RECT  6.040 -0.250 6.300 0.755 ;
        RECT  4.800 -0.250 6.040 0.250 ;
        RECT  4.200 -0.250 4.800 0.405 ;
        RECT  1.690 -0.250 4.200 0.250 ;
        RECT  1.430 -0.250 1.690 0.405 ;
        RECT  0.360 -0.250 1.430 0.250 ;
        RECT  0.360 1.035 0.385 1.295 ;
        RECT  0.125 -0.250 0.360 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.755 3.440 11.040 3.940 ;
        RECT  10.495 2.255 10.755 3.940 ;
        RECT  9.735 3.440 10.495 3.940 ;
        RECT  9.475 2.900 9.735 3.940 ;
        RECT  8.030 3.440 9.475 3.940 ;
        RECT  7.770 2.895 8.030 3.940 ;
        RECT  6.265 3.440 7.770 3.940 ;
        RECT  5.325 3.100 6.265 3.940 ;
        RECT  4.060 3.440 5.325 3.940 ;
        RECT  3.800 3.285 4.060 3.940 ;
        RECT  1.770 3.440 3.800 3.940 ;
        RECT  1.510 3.285 1.770 3.940 ;
        RECT  0.385 3.440 1.510 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.495 0.640 9.655 2.715 ;
        RECT  7.150 0.640 9.495 0.800 ;
        RECT  8.615 2.555 9.495 2.715 ;
        RECT  9.060 0.980 9.220 2.215 ;
        RECT  8.060 0.980 9.060 1.140 ;
        RECT  8.720 1.320 8.880 2.370 ;
        RECT  8.330 1.320 8.720 1.480 ;
        RECT  6.970 2.210 8.720 2.370 ;
        RECT  8.355 2.555 8.615 2.930 ;
        RECT  8.380 1.750 8.540 2.030 ;
        RECT  7.320 1.870 8.380 2.030 ;
        RECT  7.140 2.555 8.355 2.715 ;
        RECT  7.900 0.980 8.060 1.645 ;
        RECT  7.220 1.385 7.320 2.030 ;
        RECT  7.160 1.190 7.220 2.030 ;
        RECT  7.060 1.190 7.160 1.645 ;
        RECT  6.890 0.640 7.150 0.955 ;
        RECT  6.880 2.555 7.140 3.155 ;
        RECT  6.515 1.190 7.060 1.350 ;
        RECT  6.830 1.865 6.970 2.370 ;
        RECT  6.670 1.530 6.830 2.370 ;
        RECT  6.020 1.530 6.670 1.690 ;
        RECT  6.485 2.210 6.670 2.370 ;
        RECT  6.355 1.000 6.515 1.350 ;
        RECT  6.145 1.870 6.490 2.030 ;
        RECT  6.325 2.210 6.485 2.920 ;
        RECT  5.680 1.000 6.355 1.160 ;
        RECT  4.600 2.760 6.325 2.920 ;
        RECT  5.985 1.870 6.145 2.580 ;
        RECT  5.860 1.340 6.020 1.690 ;
        RECT  5.000 2.420 5.985 2.580 ;
        RECT  5.680 0.495 5.790 0.755 ;
        RECT  5.520 0.495 5.680 2.240 ;
        RECT  3.780 0.665 5.520 0.825 ;
        RECT  5.410 2.080 5.520 2.240 ;
        RECT  5.180 1.005 5.340 1.265 ;
        RECT  5.020 1.105 5.180 1.930 ;
        RECT  5.000 1.770 5.020 1.930 ;
        RECT  4.840 1.770 5.000 2.580 ;
        RECT  3.260 1.430 4.840 1.590 ;
        RECT  3.570 1.770 4.840 1.930 ;
        RECT  4.740 2.320 4.840 2.580 ;
        RECT  4.440 2.760 4.600 3.195 ;
        RECT  3.440 1.085 4.440 1.245 ;
        RECT  4.340 2.935 4.440 3.195 ;
        RECT  3.510 2.935 4.340 3.095 ;
        RECT  3.620 0.430 3.780 0.825 ;
        RECT  3.090 0.430 3.620 0.590 ;
        RECT  3.250 2.915 3.510 3.095 ;
        RECT  3.280 0.770 3.440 1.245 ;
        RECT  2.800 0.770 3.280 0.930 ;
        RECT  3.100 1.430 3.260 2.715 ;
        RECT  2.920 2.935 3.250 3.095 ;
        RECT  2.940 1.110 3.100 1.590 ;
        RECT  2.760 1.940 2.920 3.095 ;
        RECT  2.760 0.530 2.800 0.930 ;
        RECT  2.600 0.530 2.760 2.100 ;
        RECT  2.540 0.530 2.600 0.690 ;
        RECT  2.420 2.560 2.580 3.025 ;
        RECT  2.260 0.850 2.420 1.110 ;
        RECT  0.965 2.865 2.420 3.025 ;
        RECT  2.175 0.850 2.260 1.010 ;
        RECT  2.015 0.615 2.175 1.010 ;
        RECT  0.800 0.615 2.015 0.775 ;
        RECT  1.530 1.135 1.790 1.440 ;
        RECT  0.955 1.135 1.530 1.295 ;
        RECT  0.855 2.185 1.185 2.345 ;
        RECT  0.705 2.865 0.965 3.125 ;
        RECT  0.855 1.035 0.955 1.295 ;
        RECT  0.695 1.035 0.855 2.345 ;
        RECT  0.540 0.505 0.800 0.775 ;
        RECT  0.555 1.955 0.695 2.215 ;
    END
END SDFFQX4

MACRO SDFFQX2
    CLASS CORE ;
    FOREIGN SDFFQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.490 1.310 2.005 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.200 1.980 2.360 ;
        RECT  1.505 2.110 1.715 2.685 ;
        RECT  0.375 2.525 1.505 2.685 ;
        RECT  0.215 1.475 0.375 2.685 ;
        RECT  0.125 1.475 0.215 2.175 ;
        RECT  0.115 1.475 0.125 1.765 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.060 0.695 9.075 3.015 ;
        RECT  8.800 0.560 9.060 3.015 ;
        RECT  8.730 2.075 8.800 3.015 ;
        END
        ANTENNADIFFAREA     0.7272 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 1.595 2.175 1.990 ;
        RECT  1.875 1.625 1.935 1.990 ;
        RECT  1.840 1.660 1.875 1.920 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.955 2.110 4.475 2.400 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.470 -0.250 9.200 0.250 ;
        RECT  7.530 -0.250 8.470 0.405 ;
        RECT  5.710 -0.250 7.530 0.250 ;
        RECT  5.450 -0.250 5.710 0.735 ;
        RECT  4.200 -0.250 5.450 0.250 ;
        RECT  3.940 -0.250 4.200 0.405 ;
        RECT  1.690 -0.250 3.940 0.250 ;
        RECT  1.430 -0.250 1.690 0.405 ;
        RECT  0.360 -0.250 1.430 0.250 ;
        RECT  0.360 1.035 0.385 1.295 ;
        RECT  0.125 -0.250 0.360 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.480 3.440 9.200 3.940 ;
        RECT  8.220 2.855 8.480 3.940 ;
        RECT  7.490 3.440 8.220 3.940 ;
        RECT  7.230 2.875 7.490 3.940 ;
        RECT  5.845 3.440 7.230 3.940 ;
        RECT  5.245 3.285 5.845 3.940 ;
        RECT  3.940 3.440 5.245 3.940 ;
        RECT  3.680 3.285 3.940 3.940 ;
        RECT  1.875 3.440 3.680 3.940 ;
        RECT  1.615 3.285 1.875 3.940 ;
        RECT  0.385 3.440 1.615 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.510 1.495 8.560 1.755 ;
        RECT  8.350 0.590 8.510 2.675 ;
        RECT  7.370 0.590 8.350 0.750 ;
        RECT  8.300 1.495 8.350 1.755 ;
        RECT  6.820 2.515 8.350 2.675 ;
        RECT  7.975 1.035 8.150 1.295 ;
        RECT  7.975 2.075 8.075 2.335 ;
        RECT  7.890 1.035 7.975 2.335 ;
        RECT  7.815 1.085 7.890 2.335 ;
        RECT  7.440 1.435 7.815 1.645 ;
        RECT  7.180 1.385 7.440 1.645 ;
        RECT  7.210 0.525 7.370 0.750 ;
        RECT  6.460 0.525 7.210 0.685 ;
        RECT  6.980 0.905 7.030 1.165 ;
        RECT  6.820 0.905 6.980 1.865 ;
        RECT  6.770 0.905 6.820 1.165 ;
        RECT  6.650 1.705 6.820 1.865 ;
        RECT  6.560 2.515 6.820 3.115 ;
        RECT  6.210 0.905 6.770 1.065 ;
        RECT  6.550 1.705 6.650 1.965 ;
        RECT  6.155 1.275 6.550 1.435 ;
        RECT  6.390 1.705 6.550 2.300 ;
        RECT  6.190 2.140 6.390 2.300 ;
        RECT  6.050 0.905 6.210 1.095 ;
        RECT  6.030 2.140 6.190 3.095 ;
        RECT  5.845 1.755 6.170 1.915 ;
        RECT  5.995 1.275 6.155 1.570 ;
        RECT  5.590 0.935 6.050 1.095 ;
        RECT  4.490 2.935 6.030 3.095 ;
        RECT  5.250 1.410 5.995 1.570 ;
        RECT  5.685 1.755 5.845 2.685 ;
        RECT  4.910 2.525 5.685 2.685 ;
        RECT  5.430 0.935 5.590 1.195 ;
        RECT  5.250 2.075 5.465 2.335 ;
        RECT  5.205 0.675 5.250 2.335 ;
        RECT  5.140 0.675 5.205 2.285 ;
        RECT  5.090 0.495 5.140 2.285 ;
        RECT  4.880 0.495 5.090 0.835 ;
        RECT  4.750 1.055 4.910 2.685 ;
        RECT  3.755 0.675 4.880 0.835 ;
        RECT  4.520 1.055 4.750 1.215 ;
        RECT  3.590 1.770 4.750 1.930 ;
        RECT  4.680 2.425 4.750 2.685 ;
        RECT  3.150 1.430 4.570 1.590 ;
        RECT  4.230 2.935 4.490 3.195 ;
        RECT  3.400 2.935 4.230 3.100 ;
        RECT  3.205 1.080 4.200 1.240 ;
        RECT  3.595 0.430 3.755 0.835 ;
        RECT  3.020 0.430 3.595 0.590 ;
        RECT  3.330 1.770 3.590 2.030 ;
        RECT  3.140 2.915 3.400 3.100 ;
        RECT  3.045 0.770 3.205 1.240 ;
        RECT  2.990 1.430 3.150 2.720 ;
        RECT  2.810 2.940 3.140 3.100 ;
        RECT  2.770 0.770 3.045 0.930 ;
        RECT  2.860 1.430 2.990 1.590 ;
        RECT  2.700 1.110 2.860 1.590 ;
        RECT  2.650 1.940 2.810 3.100 ;
        RECT  2.515 0.655 2.770 0.930 ;
        RECT  2.515 1.940 2.650 2.100 ;
        RECT  2.510 0.655 2.515 2.100 ;
        RECT  2.355 0.770 2.510 2.100 ;
        RECT  2.370 3.100 2.470 3.260 ;
        RECT  2.210 2.865 2.370 3.260 ;
        RECT  2.175 0.430 2.330 0.590 ;
        RECT  0.965 2.865 2.210 3.025 ;
        RECT  2.015 0.430 2.175 0.775 ;
        RECT  0.800 0.615 2.015 0.775 ;
        RECT  1.530 1.135 1.790 1.440 ;
        RECT  0.955 1.135 1.530 1.295 ;
        RECT  0.855 2.185 1.185 2.345 ;
        RECT  0.705 2.865 0.965 3.125 ;
        RECT  0.855 1.035 0.955 1.295 ;
        RECT  0.695 1.035 0.855 2.345 ;
        RECT  0.540 0.455 0.800 0.775 ;
        RECT  0.555 1.955 0.695 2.215 ;
    END
END SDFFQX2

MACRO SDFFQX1
    CLASS CORE ;
    FOREIGN SDFFQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.490 1.310 2.005 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.170 1.980 2.430 ;
        RECT  1.505 2.110 1.715 2.765 ;
        RECT  0.375 2.605 1.505 2.765 ;
        RECT  0.215 1.475 0.375 2.765 ;
        RECT  0.125 1.475 0.215 2.175 ;
        RECT  0.115 1.475 0.125 1.765 ;
        END
        ANTENNAGATEAREA     0.0897 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.465 0.600 8.625 2.755 ;
        RECT  8.430 0.600 8.465 0.760 ;
        RECT  8.195 2.595 8.465 2.755 ;
        RECT  8.155 0.495 8.430 0.760 ;
        RECT  7.935 2.595 8.195 3.195 ;
        RECT  7.945 0.470 8.155 0.760 ;
        END
        ANTENNADIFFAREA     0.3366 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 1.595 2.175 1.990 ;
        RECT  1.875 1.625 1.935 1.990 ;
        RECT  1.840 1.670 1.875 1.930 ;
        END
        ANTENNAGATEAREA     0.0403 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 2.110 4.595 2.400 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.705 -0.250 8.740 0.250 ;
        RECT  7.445 -0.250 7.705 0.595 ;
        RECT  6.035 -0.250 7.445 0.250 ;
        RECT  5.775 -0.250 6.035 0.945 ;
        RECT  4.440 -0.250 5.775 0.250 ;
        RECT  3.840 -0.250 4.440 0.625 ;
        RECT  1.690 -0.250 3.840 0.250 ;
        RECT  1.430 -0.250 1.690 0.405 ;
        RECT  0.360 -0.250 1.430 0.250 ;
        RECT  0.360 1.035 0.385 1.295 ;
        RECT  0.125 -0.250 0.360 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.645 3.440 8.740 3.940 ;
        RECT  7.385 2.500 7.645 3.940 ;
        RECT  5.860 3.440 7.385 3.940 ;
        RECT  5.600 3.285 5.860 3.940 ;
        RECT  4.850 3.440 5.600 3.940 ;
        RECT  4.590 3.285 4.850 3.940 ;
        RECT  3.940 3.440 4.590 3.940 ;
        RECT  3.680 3.285 3.940 3.940 ;
        RECT  1.875 3.440 3.680 3.940 ;
        RECT  1.615 3.285 1.875 3.940 ;
        RECT  0.385 3.440 1.615 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.235 1.035 8.285 1.295 ;
        RECT  8.075 1.035 8.235 2.320 ;
        RECT  8.025 1.035 8.075 1.295 ;
        RECT  7.975 2.055 8.075 2.320 ;
        RECT  7.400 2.055 7.975 2.215 ;
        RECT  7.800 1.495 7.865 1.755 ;
        RECT  7.640 1.240 7.800 1.755 ;
        RECT  6.940 1.240 7.640 1.400 ;
        RECT  7.240 1.590 7.400 2.215 ;
        RECT  7.140 1.590 7.240 1.850 ;
        RECT  6.855 0.435 7.115 0.695 ;
        RECT  6.935 0.875 6.940 1.400 ;
        RECT  6.775 0.875 6.935 2.765 ;
        RECT  6.405 0.535 6.855 0.695 ;
        RECT  6.595 0.875 6.775 1.035 ;
        RECT  6.720 2.605 6.775 2.765 ;
        RECT  6.460 2.605 6.720 2.865 ;
        RECT  6.455 2.040 6.595 2.300 ;
        RECT  6.405 1.305 6.455 2.300 ;
        RECT  6.295 0.535 6.405 2.300 ;
        RECT  6.245 0.535 6.295 1.465 ;
        RECT  6.190 2.140 6.295 2.300 ;
        RECT  5.845 1.305 6.245 1.465 ;
        RECT  6.030 2.140 6.190 3.105 ;
        RECT  5.855 1.685 6.115 1.945 ;
        RECT  4.450 2.945 6.030 3.105 ;
        RECT  5.845 1.785 5.855 1.945 ;
        RECT  5.685 1.205 5.845 1.465 ;
        RECT  5.685 1.785 5.845 2.750 ;
        RECT  4.980 2.590 5.685 2.750 ;
        RECT  5.345 0.430 5.505 2.290 ;
        RECT  5.120 0.430 5.345 0.805 ;
        RECT  5.170 2.030 5.345 2.290 ;
        RECT  5.005 1.070 5.165 1.335 ;
        RECT  4.745 0.430 5.120 0.590 ;
        RECT  4.980 1.175 5.005 1.335 ;
        RECT  4.820 1.175 4.980 2.750 ;
        RECT  3.730 1.770 4.820 1.930 ;
        RECT  3.150 1.430 4.505 1.590 ;
        RECT  4.190 2.580 4.450 3.105 ;
        RECT  4.015 0.935 4.275 1.195 ;
        RECT  3.400 2.940 4.190 3.105 ;
        RECT  3.490 1.035 4.015 1.195 ;
        RECT  3.630 1.770 3.730 1.935 ;
        RECT  3.370 1.770 3.630 2.030 ;
        RECT  3.330 0.770 3.490 1.195 ;
        RECT  3.140 2.915 3.400 3.105 ;
        RECT  2.560 0.770 3.330 0.930 ;
        RECT  2.990 1.430 3.150 2.660 ;
        RECT  2.810 2.945 3.140 3.105 ;
        RECT  2.900 1.430 2.990 1.590 ;
        RECT  2.740 1.110 2.900 1.590 ;
        RECT  2.650 1.940 2.810 3.105 ;
        RECT  2.560 1.940 2.650 2.100 ;
        RECT  2.400 0.770 2.560 2.100 ;
        RECT  2.310 2.945 2.470 3.245 ;
        RECT  2.370 1.305 2.400 1.565 ;
        RECT  2.220 0.430 2.330 0.590 ;
        RECT  0.965 2.945 2.310 3.105 ;
        RECT  2.060 0.430 2.220 0.775 ;
        RECT  0.800 0.615 2.060 0.775 ;
        RECT  1.530 1.135 1.790 1.440 ;
        RECT  0.955 1.135 1.530 1.295 ;
        RECT  0.855 2.265 1.185 2.425 ;
        RECT  0.705 2.945 0.965 3.205 ;
        RECT  0.855 1.035 0.955 1.295 ;
        RECT  0.695 1.035 0.855 2.425 ;
        RECT  0.540 0.505 0.800 0.775 ;
        RECT  0.555 1.955 0.695 2.215 ;
    END
END SDFFQX1

MACRO SDFFX4
    CLASS CORE ;
    FOREIGN SDFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.340 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.505 1.405 1.895 ;
        RECT  1.045 1.505 1.255 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.065 1.975 2.325 ;
        RECT  1.665 2.110 1.715 2.400 ;
        RECT  1.505 2.110 1.665 2.670 ;
        RECT  0.350 2.510 1.505 2.670 ;
        RECT  0.350 1.480 0.445 1.740 ;
        RECT  0.190 1.480 0.350 2.670 ;
        RECT  0.185 1.480 0.190 2.175 ;
        RECT  0.125 1.700 0.185 2.175 ;
        END
        ANTENNAGATEAREA     0.1352 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.685 1.035 12.755 2.585 ;
        RECT  12.495 0.695 12.685 2.895 ;
        RECT  12.425 0.695 12.495 1.295 ;
        RECT  12.425 1.955 12.495 2.895 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.665 1.515 11.835 1.765 ;
        RECT  11.405 0.695 11.665 2.215 ;
        RECT  11.165 1.290 11.405 1.990 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.700 2.635 2.165 ;
        RECT  2.195 1.755 2.425 2.165 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.525 1.810 4.785 2.070 ;
        RECT  4.475 1.910 4.525 2.070 ;
        RECT  4.315 1.910 4.475 2.400 ;
        RECT  4.265 2.110 4.315 2.400 ;
        END
        ANTENNAGATEAREA     0.2002 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.195 -0.250 13.340 0.250 ;
        RECT  12.935 -0.250 13.195 1.095 ;
        RECT  12.175 -0.250 12.935 0.250 ;
        RECT  11.915 -0.250 12.175 1.095 ;
        RECT  11.155 -0.250 11.915 0.250 ;
        RECT  10.895 -0.250 11.155 0.755 ;
        RECT  10.240 -0.250 10.895 0.250 ;
        RECT  9.995 -0.250 10.240 1.250 ;
        RECT  9.925 -0.250 9.995 0.405 ;
        RECT  8.365 -0.250 9.925 0.250 ;
        RECT  8.105 -0.250 8.365 0.575 ;
        RECT  6.695 -0.250 8.105 0.250 ;
        RECT  6.435 -0.250 6.695 0.895 ;
        RECT  5.005 -0.250 6.435 0.250 ;
        RECT  4.745 -0.250 5.005 0.745 ;
        RECT  4.095 -0.250 4.745 0.250 ;
        RECT  3.835 -0.250 4.095 0.945 ;
        RECT  1.785 -0.250 3.835 0.250 ;
        RECT  1.525 -0.250 1.785 0.405 ;
        RECT  0.385 -0.250 1.525 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.195 3.440 13.340 3.940 ;
        RECT  12.935 2.255 13.195 3.940 ;
        RECT  12.175 3.440 12.935 3.940 ;
        RECT  11.915 2.935 12.175 3.940 ;
        RECT  11.155 3.440 11.915 3.940 ;
        RECT  10.895 2.935 11.155 3.940 ;
        RECT  10.215 3.440 10.895 3.940 ;
        RECT  9.955 2.410 10.215 3.940 ;
        RECT  8.365 3.440 9.955 3.940 ;
        RECT  8.105 2.715 8.365 3.940 ;
        RECT  6.665 3.440 8.105 3.940 ;
        RECT  6.405 3.285 6.665 3.940 ;
        RECT  5.165 3.440 6.405 3.940 ;
        RECT  4.905 3.285 5.165 3.940 ;
        RECT  4.105 3.440 4.905 3.940 ;
        RECT  3.845 3.285 4.105 3.940 ;
        RECT  1.875 3.440 3.845 3.940 ;
        RECT  1.615 3.285 1.875 3.940 ;
        RECT  0.385 3.440 1.615 3.940 ;
        RECT  0.125 2.870 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.215 1.515 12.315 1.775 ;
        RECT  12.055 1.515 12.215 2.585 ;
        RECT  10.755 2.425 12.055 2.585 ;
        RECT  10.705 1.035 10.755 1.295 ;
        RECT  10.705 1.985 10.755 2.585 ;
        RECT  10.545 1.035 10.705 2.585 ;
        RECT  10.495 1.035 10.545 1.295 ;
        RECT  10.495 1.985 10.545 2.585 ;
        RECT  9.730 1.985 10.495 2.145 ;
        RECT  10.105 1.515 10.365 1.775 ;
        RECT  9.815 1.565 10.105 1.775 ;
        RECT  9.655 0.755 9.815 1.775 ;
        RECT  9.730 2.855 9.775 3.115 ;
        RECT  9.570 1.985 9.730 3.115 ;
        RECT  9.215 0.755 9.655 0.915 ;
        RECT  9.390 1.615 9.655 1.775 ;
        RECT  9.515 2.855 9.570 3.115 ;
        RECT  9.045 1.145 9.475 1.405 ;
        RECT  9.230 1.615 9.390 2.535 ;
        RECT  9.215 2.375 9.230 2.535 ;
        RECT  8.955 0.705 9.215 0.965 ;
        RECT  8.955 2.375 9.215 2.990 ;
        RECT  8.885 1.145 9.045 2.195 ;
        RECT  7.255 0.755 8.955 0.915 ;
        RECT  7.515 2.375 8.955 2.535 ;
        RECT  8.510 1.145 8.885 1.305 ;
        RECT  8.785 1.805 8.885 2.195 ;
        RECT  7.205 1.805 8.785 1.965 ;
        RECT  8.350 1.095 8.510 1.305 ;
        RECT  6.525 1.095 8.350 1.255 ;
        RECT  6.865 1.435 8.165 1.595 ;
        RECT  7.255 2.375 7.515 2.975 ;
        RECT  7.045 1.805 7.205 2.170 ;
        RECT  6.755 2.010 7.045 2.170 ;
        RECT  6.705 1.435 6.865 1.830 ;
        RECT  6.595 2.010 6.755 3.105 ;
        RECT  6.375 1.670 6.705 1.830 ;
        RECT  3.565 2.945 6.595 3.105 ;
        RECT  6.365 1.095 6.525 1.390 ;
        RECT  6.215 1.670 6.375 2.765 ;
        RECT  6.355 1.230 6.365 1.390 ;
        RECT  6.095 1.230 6.355 1.490 ;
        RECT  5.515 2.605 6.215 2.765 ;
        RECT  5.915 0.790 6.185 1.050 ;
        RECT  5.915 2.045 5.965 2.305 ;
        RECT  5.755 0.470 5.915 2.305 ;
        RECT  5.565 0.470 5.755 0.630 ;
        RECT  5.705 2.045 5.755 2.305 ;
        RECT  5.515 0.825 5.565 1.085 ;
        RECT  5.355 0.825 5.515 2.765 ;
        RECT  5.305 0.825 5.355 1.085 ;
        RECT  4.045 2.605 5.355 2.765 ;
        RECT  4.900 1.265 5.160 1.630 ;
        RECT  3.315 1.470 4.900 1.630 ;
        RECT  4.345 0.995 4.605 1.285 ;
        RECT  3.655 1.125 4.345 1.285 ;
        RECT  3.885 1.915 4.045 2.765 ;
        RECT  3.785 1.915 3.885 2.175 ;
        RECT  3.495 0.545 3.655 1.285 ;
        RECT  3.305 2.895 3.565 3.155 ;
        RECT  2.825 0.545 3.495 0.705 ;
        RECT  3.165 0.985 3.315 2.695 ;
        RECT  2.975 2.945 3.305 3.105 ;
        RECT  3.155 0.885 3.165 2.695 ;
        RECT  3.005 0.885 3.155 1.145 ;
        RECT  2.825 1.325 2.975 3.105 ;
        RECT  2.815 0.545 2.825 3.105 ;
        RECT  2.665 0.545 2.815 1.485 ;
        RECT  2.615 1.325 2.665 1.485 ;
        RECT  2.525 2.540 2.625 2.800 ;
        RECT  2.365 2.540 2.525 3.010 ;
        RECT  2.325 0.585 2.485 1.145 ;
        RECT  0.985 2.850 2.365 3.010 ;
        RECT  1.010 0.585 2.325 0.745 ;
        RECT  1.785 1.320 1.885 1.580 ;
        RECT  1.625 1.135 1.785 1.580 ;
        RECT  0.815 1.135 1.625 1.295 ;
        RECT  0.815 2.170 1.185 2.330 ;
        RECT  0.850 0.470 1.010 0.745 ;
        RECT  0.725 2.850 0.985 3.110 ;
        RECT  0.635 0.470 0.850 0.630 ;
        RECT  0.785 1.035 0.815 1.295 ;
        RECT  0.785 2.070 0.815 2.330 ;
        RECT  0.625 1.035 0.785 2.330 ;
        RECT  0.555 1.035 0.625 1.295 ;
        RECT  0.555 2.070 0.625 2.330 ;
    END
END SDFFX4

MACRO SDFFX2
    CLASS CORE ;
    FOREIGN SDFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.475 1.310 1.735 ;
        RECT  1.255 1.475 1.260 1.925 ;
        RECT  1.050 1.475 1.255 1.990 ;
        RECT  1.045 1.700 1.050 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.170 1.980 2.430 ;
        RECT  1.505 2.110 1.715 2.765 ;
        RECT  0.325 2.605 1.505 2.765 ;
        RECT  0.335 1.575 0.375 1.835 ;
        RECT  0.325 1.575 0.335 2.175 ;
        RECT  0.165 1.575 0.325 2.765 ;
        RECT  0.115 1.575 0.165 2.175 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.245 0.695 10.455 3.045 ;
        RECT  10.195 0.695 10.245 1.295 ;
        RECT  10.195 2.105 10.245 3.045 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.900 1.700 9.075 1.990 ;
        RECT  8.865 0.495 9.055 0.755 ;
        RECT  8.770 1.700 8.900 2.215 ;
        RECT  8.795 0.495 8.865 0.760 ;
        RECT  8.770 0.595 8.795 0.760 ;
        RECT  8.610 0.595 8.770 2.215 ;
        END
        ANTENNADIFFAREA     0.6173 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.670 2.305 1.990 ;
        RECT  1.840 1.670 1.965 1.930 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 2.110 4.595 2.400 ;
        END
        ANTENNAGATEAREA     0.1144 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.915 -0.250 10.580 0.250 ;
        RECT  9.655 -0.250 9.915 0.645 ;
        RECT  8.510 -0.250 9.655 0.250 ;
        RECT  8.250 -0.250 8.510 0.405 ;
        RECT  6.360 -0.250 8.250 0.250 ;
        RECT  6.100 -0.250 6.360 0.635 ;
        RECT  4.960 -0.250 6.100 0.250 ;
        RECT  4.020 -0.250 4.960 0.405 ;
        RECT  1.690 -0.250 4.020 0.250 ;
        RECT  1.430 -0.250 1.690 0.405 ;
        RECT  0.360 -0.250 1.430 0.250 ;
        RECT  0.360 1.035 0.385 1.295 ;
        RECT  0.125 -0.250 0.360 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.915 3.440 10.580 3.940 ;
        RECT  9.655 2.205 9.915 3.940 ;
        RECT  8.350 3.440 9.655 3.940 ;
        RECT  8.090 2.890 8.350 3.940 ;
        RECT  6.160 3.440 8.090 3.940 ;
        RECT  5.900 3.285 6.160 3.940 ;
        RECT  5.140 3.440 5.900 3.940 ;
        RECT  4.880 3.285 5.140 3.940 ;
        RECT  4.080 3.440 4.880 3.940 ;
        RECT  3.820 3.285 4.080 3.940 ;
        RECT  1.875 3.440 3.820 3.940 ;
        RECT  1.615 3.285 1.875 3.940 ;
        RECT  0.385 3.440 1.615 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.455 1.585 10.055 1.845 ;
        RECT  9.295 1.035 9.455 2.725 ;
        RECT  9.195 1.035 9.295 1.295 ;
        RECT  9.105 2.465 9.295 2.725 ;
        RECT  7.910 2.465 9.105 2.625 ;
        RECT  8.180 0.610 8.340 2.130 ;
        RECT  8.070 0.610 8.180 0.770 ;
        RECT  7.565 1.970 8.180 2.130 ;
        RECT  7.910 0.470 8.070 0.770 ;
        RECT  7.780 0.950 7.940 1.790 ;
        RECT  7.290 0.470 7.910 0.630 ;
        RECT  7.750 2.465 7.910 2.905 ;
        RECT  7.730 0.950 7.780 1.110 ;
        RECT  7.225 1.630 7.780 1.790 ;
        RECT  7.650 2.645 7.750 2.905 ;
        RECT  7.520 0.810 7.730 1.110 ;
        RECT  6.860 1.290 7.600 1.450 ;
        RECT  7.405 1.970 7.565 2.455 ;
        RECT  7.470 0.810 7.520 1.075 ;
        RECT  6.170 0.915 7.470 1.075 ;
        RECT  7.015 2.295 7.405 2.455 ;
        RECT  7.130 0.470 7.290 0.735 ;
        RECT  7.065 1.630 7.225 2.115 ;
        RECT  6.510 1.955 7.065 2.115 ;
        RECT  6.755 2.295 7.015 2.895 ;
        RECT  6.700 1.275 6.860 1.450 ;
        RECT  5.830 1.275 6.700 1.435 ;
        RECT  6.350 1.955 6.510 3.105 ;
        RECT  4.590 2.945 6.350 3.105 ;
        RECT  6.170 1.615 6.270 1.775 ;
        RECT  6.010 0.815 6.170 1.075 ;
        RECT  6.010 1.615 6.170 2.735 ;
        RECT  5.080 2.575 6.010 2.735 ;
        RECT  5.670 0.595 5.830 2.225 ;
        RECT  5.540 0.595 5.670 0.755 ;
        RECT  5.570 2.015 5.670 2.225 ;
        RECT  5.310 2.015 5.570 2.275 ;
        RECT  5.280 0.495 5.540 0.755 ;
        RECT  5.330 1.015 5.490 1.645 ;
        RECT  5.080 1.485 5.330 1.645 ;
        RECT  3.780 0.595 5.280 0.755 ;
        RECT  4.920 1.485 5.080 2.735 ;
        RECT  3.830 1.770 4.920 1.930 ;
        RECT  3.290 1.430 4.740 1.590 ;
        RECT  3.440 1.060 4.600 1.220 ;
        RECT  4.330 2.595 4.590 3.105 ;
        RECT  3.540 2.945 4.330 3.105 ;
        RECT  3.570 1.770 3.830 2.030 ;
        RECT  3.620 0.470 3.780 0.755 ;
        RECT  3.280 2.915 3.540 3.175 ;
        RECT  3.280 0.670 3.440 1.220 ;
        RECT  3.130 1.430 3.290 2.650 ;
        RECT  2.760 0.670 3.280 0.830 ;
        RECT  2.950 2.915 3.280 3.075 ;
        RECT  3.100 1.430 3.130 1.590 ;
        RECT  2.940 1.010 3.100 1.590 ;
        RECT  2.790 1.940 2.950 3.075 ;
        RECT  2.760 1.940 2.790 2.100 ;
        RECT  2.600 0.670 2.760 2.100 ;
        RECT  2.450 2.390 2.610 3.105 ;
        RECT  2.500 1.375 2.600 1.635 ;
        RECT  0.965 2.945 2.450 3.105 ;
        RECT  2.260 0.615 2.420 1.195 ;
        RECT  0.800 0.615 2.260 0.775 ;
        RECT  1.530 1.135 1.790 1.425 ;
        RECT  0.955 1.135 1.530 1.295 ;
        RECT  0.855 2.265 1.185 2.425 ;
        RECT  0.705 2.945 0.965 3.205 ;
        RECT  0.855 1.035 0.955 1.295 ;
        RECT  0.695 1.035 0.855 2.425 ;
        RECT  0.590 0.505 0.800 0.775 ;
        RECT  0.555 1.955 0.695 2.215 ;
        RECT  0.540 0.505 0.590 0.665 ;
    END
END SDFFX2

MACRO SDFFX1
    CLASS CORE ;
    FOREIGN SDFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.475 1.310 1.735 ;
        RECT  1.255 1.475 1.260 1.925 ;
        RECT  1.050 1.475 1.255 1.990 ;
        RECT  1.045 1.700 1.050 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.170 1.980 2.430 ;
        RECT  1.505 2.110 1.715 2.765 ;
        RECT  0.375 2.605 1.505 2.765 ;
        RECT  0.375 1.505 0.500 1.765 ;
        RECT  0.215 1.505 0.375 2.765 ;
        RECT  0.125 1.925 0.215 2.335 ;
        END
        ANTENNAGATEAREA     0.0923 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.520 1.100 9.535 2.715 ;
        RECT  9.325 1.030 9.520 2.715 ;
        RECT  9.260 1.030 9.325 1.290 ;
        RECT  9.260 2.115 9.325 2.715 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.075 0.945 9.080 2.665 ;
        RECT  9.025 0.880 9.075 2.665 ;
        RECT  8.920 0.715 9.025 2.665 ;
        RECT  8.865 0.715 8.920 1.170 ;
        RECT  8.865 2.335 8.920 2.665 ;
        RECT  8.400 0.715 8.865 0.875 ;
        RECT  8.460 2.505 8.865 2.665 ;
        RECT  8.200 2.505 8.460 3.195 ;
        RECT  8.140 0.615 8.400 0.875 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.670 2.305 1.990 ;
        RECT  1.840 1.670 1.965 1.930 ;
        END
        ANTENNAGATEAREA     0.0429 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 2.110 4.595 2.400 ;
        END
        ANTENNAGATEAREA     0.0793 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.000 -0.250 9.660 0.250 ;
        RECT  8.740 -0.250 9.000 0.405 ;
        RECT  7.850 -0.250 8.740 0.250 ;
        RECT  7.590 -0.250 7.850 0.405 ;
        RECT  6.170 -0.250 7.590 0.250 ;
        RECT  5.910 -0.250 6.170 0.945 ;
        RECT  4.720 -0.250 5.910 0.250 ;
        RECT  3.780 -0.250 4.720 0.625 ;
        RECT  1.690 -0.250 3.780 0.250 ;
        RECT  1.430 -0.250 1.690 0.405 ;
        RECT  0.360 -0.250 1.430 0.250 ;
        RECT  0.360 1.035 0.385 1.295 ;
        RECT  0.125 -0.250 0.360 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.970 3.440 9.660 3.940 ;
        RECT  8.710 2.875 8.970 3.940 ;
        RECT  7.920 3.440 8.710 3.940 ;
        RECT  7.660 2.875 7.920 3.940 ;
        RECT  6.000 3.440 7.660 3.940 ;
        RECT  5.740 3.285 6.000 3.940 ;
        RECT  5.140 3.440 5.740 3.940 ;
        RECT  4.880 3.285 5.140 3.940 ;
        RECT  4.080 3.440 4.880 3.940 ;
        RECT  3.820 3.285 4.080 3.940 ;
        RECT  1.875 3.440 3.820 3.940 ;
        RECT  1.615 3.285 1.875 3.940 ;
        RECT  0.385 3.440 1.615 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.490 1.625 8.740 1.885 ;
        RECT  8.460 1.125 8.490 2.275 ;
        RECT  8.330 1.125 8.460 2.325 ;
        RECT  8.230 1.125 8.330 1.385 ;
        RECT  8.200 2.065 8.330 2.325 ;
        RECT  7.670 2.065 8.200 2.225 ;
        RECT  8.050 1.565 8.150 1.825 ;
        RECT  7.890 1.240 8.050 1.825 ;
        RECT  7.230 1.240 7.890 1.400 ;
        RECT  7.510 1.695 7.670 2.225 ;
        RECT  7.410 1.695 7.510 1.955 ;
        RECT  6.540 0.555 7.310 0.715 ;
        RECT  7.070 0.895 7.230 2.580 ;
        RECT  6.820 0.895 7.070 1.155 ;
        RECT  6.980 2.420 7.070 2.580 ;
        RECT  6.720 2.420 6.980 3.020 ;
        RECT  6.540 1.945 6.880 2.205 ;
        RECT  6.380 0.555 6.540 3.075 ;
        RECT  6.040 1.305 6.380 1.465 ;
        RECT  4.590 2.915 6.380 3.075 ;
        RECT  6.040 1.685 6.200 2.735 ;
        RECT  5.880 1.205 6.040 1.465 ;
        RECT  4.980 2.575 6.040 2.735 ;
        RECT  5.570 0.460 5.700 2.160 ;
        RECT  5.540 0.460 5.570 2.275 ;
        RECT  5.310 0.460 5.540 0.815 ;
        RECT  5.310 2.000 5.540 2.275 ;
        RECT  5.200 1.065 5.360 1.325 ;
        RECT  4.940 0.460 5.310 0.620 ;
        RECT  4.980 1.165 5.200 1.325 ;
        RECT  4.820 1.165 4.980 2.735 ;
        RECT  3.830 1.770 4.820 1.930 ;
        RECT  3.290 1.430 4.640 1.590 ;
        RECT  4.330 2.595 4.590 3.075 ;
        RECT  4.210 0.935 4.470 1.195 ;
        RECT  3.540 2.915 4.330 3.075 ;
        RECT  3.490 0.935 4.210 1.095 ;
        RECT  3.570 1.770 3.830 2.030 ;
        RECT  3.280 2.865 3.540 3.125 ;
        RECT  3.330 0.585 3.490 1.095 ;
        RECT  2.760 0.585 3.330 0.745 ;
        RECT  3.130 1.430 3.290 2.650 ;
        RECT  2.950 2.915 3.280 3.075 ;
        RECT  3.100 1.430 3.130 1.590 ;
        RECT  2.940 0.935 3.100 1.590 ;
        RECT  2.790 1.940 2.950 3.075 ;
        RECT  2.760 1.940 2.790 2.100 ;
        RECT  2.600 0.585 2.760 2.100 ;
        RECT  2.450 2.430 2.610 3.105 ;
        RECT  2.500 1.375 2.600 1.635 ;
        RECT  0.965 2.945 2.450 3.105 ;
        RECT  2.260 0.615 2.420 1.195 ;
        RECT  0.800 0.615 2.260 0.775 ;
        RECT  1.530 1.135 1.790 1.425 ;
        RECT  0.955 1.135 1.530 1.295 ;
        RECT  0.855 2.265 1.185 2.425 ;
        RECT  0.705 2.945 0.965 3.205 ;
        RECT  0.855 1.035 0.955 1.295 ;
        RECT  0.695 1.035 0.855 2.425 ;
        RECT  0.540 0.455 0.800 0.775 ;
        RECT  0.555 1.955 0.695 2.215 ;
    END
END SDFFX1

MACRO SDFFXL
    CLASS CORE ;
    FOREIGN SDFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.475 1.310 1.735 ;
        RECT  1.255 1.475 1.260 1.925 ;
        RECT  1.050 1.475 1.255 1.990 ;
        RECT  1.045 1.700 1.050 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.170 1.980 2.430 ;
        RECT  1.505 2.110 1.715 2.765 ;
        RECT  0.325 2.605 1.505 2.765 ;
        RECT  0.335 1.475 0.375 1.735 ;
        RECT  0.325 1.475 0.335 2.175 ;
        RECT  0.165 1.475 0.325 2.765 ;
        RECT  0.115 1.475 0.165 2.175 ;
        END
        ANTENNAGATEAREA     0.0923 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.520 1.105 9.535 2.175 ;
        RECT  9.325 1.030 9.520 2.375 ;
        RECT  9.260 1.030 9.325 1.290 ;
        RECT  9.260 2.115 9.325 2.375 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.075 0.945 9.080 2.665 ;
        RECT  9.025 0.880 9.075 2.665 ;
        RECT  8.920 0.615 9.025 2.665 ;
        RECT  8.865 0.615 8.920 1.170 ;
        RECT  8.830 2.335 8.920 2.665 ;
        RECT  8.435 0.615 8.865 0.775 ;
        RECT  8.460 2.505 8.830 2.665 ;
        RECT  8.300 2.505 8.460 3.005 ;
        RECT  8.175 0.515 8.435 0.775 ;
        RECT  8.200 2.745 8.300 3.005 ;
        END
        ANTENNADIFFAREA     0.2221 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.670 2.305 1.990 ;
        RECT  1.840 1.670 1.965 1.930 ;
        END
        ANTENNAGATEAREA     0.0429 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 2.110 4.595 2.400 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.965 -0.250 9.660 0.250 ;
        RECT  8.705 -0.250 8.965 0.405 ;
        RECT  7.850 -0.250 8.705 0.250 ;
        RECT  7.590 -0.250 7.850 0.405 ;
        RECT  6.170 -0.250 7.590 0.250 ;
        RECT  5.910 -0.250 6.170 0.945 ;
        RECT  4.720 -0.250 5.910 0.250 ;
        RECT  3.780 -0.250 4.720 0.625 ;
        RECT  1.690 -0.250 3.780 0.250 ;
        RECT  1.430 -0.250 1.690 0.405 ;
        RECT  0.360 -0.250 1.430 0.250 ;
        RECT  0.360 1.035 0.385 1.295 ;
        RECT  0.125 -0.250 0.360 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.970 3.440 9.660 3.940 ;
        RECT  8.710 2.875 8.970 3.940 ;
        RECT  7.920 3.440 8.710 3.940 ;
        RECT  7.660 2.555 7.920 3.940 ;
        RECT  6.030 3.440 7.660 3.940 ;
        RECT  5.770 3.285 6.030 3.940 ;
        RECT  5.170 3.440 5.770 3.940 ;
        RECT  4.910 3.285 5.170 3.940 ;
        RECT  4.080 3.440 4.910 3.940 ;
        RECT  3.820 3.285 4.080 3.940 ;
        RECT  1.875 3.440 3.820 3.940 ;
        RECT  1.615 3.285 1.875 3.940 ;
        RECT  0.385 3.440 1.615 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.490 1.625 8.740 1.885 ;
        RECT  8.330 1.025 8.490 2.325 ;
        RECT  8.190 1.025 8.330 1.285 ;
        RECT  8.230 2.065 8.330 2.325 ;
        RECT  7.670 2.065 8.230 2.225 ;
        RECT  8.010 1.565 8.150 1.825 ;
        RECT  7.850 1.240 8.010 1.825 ;
        RECT  7.230 1.240 7.850 1.400 ;
        RECT  7.510 1.695 7.670 2.225 ;
        RECT  7.410 1.695 7.510 1.955 ;
        RECT  6.570 0.555 7.310 0.715 ;
        RECT  7.070 0.895 7.230 2.620 ;
        RECT  6.820 0.895 7.070 1.155 ;
        RECT  6.960 2.460 7.070 2.620 ;
        RECT  6.700 2.460 6.960 2.720 ;
        RECT  6.570 1.945 6.880 2.280 ;
        RECT  6.520 0.555 6.570 2.280 ;
        RECT  6.410 0.555 6.520 3.105 ;
        RECT  6.040 1.305 6.410 1.465 ;
        RECT  6.360 2.120 6.410 3.105 ;
        RECT  4.590 2.945 6.360 3.105 ;
        RECT  6.170 1.675 6.230 1.935 ;
        RECT  6.010 1.675 6.170 2.765 ;
        RECT  5.880 1.195 6.040 1.465 ;
        RECT  4.980 2.605 6.010 2.765 ;
        RECT  5.540 0.460 5.700 2.305 ;
        RECT  5.310 0.460 5.540 0.795 ;
        RECT  5.340 2.045 5.540 2.305 ;
        RECT  5.200 1.045 5.360 1.325 ;
        RECT  4.940 0.460 5.310 0.620 ;
        RECT  4.980 1.165 5.200 1.325 ;
        RECT  4.820 1.165 4.980 2.765 ;
        RECT  3.830 1.770 4.820 1.930 ;
        RECT  3.290 1.430 4.640 1.590 ;
        RECT  4.330 2.595 4.590 3.105 ;
        RECT  4.210 0.935 4.470 1.195 ;
        RECT  3.540 2.945 4.330 3.105 ;
        RECT  3.490 0.935 4.210 1.095 ;
        RECT  3.570 1.770 3.830 2.030 ;
        RECT  3.280 2.900 3.540 3.160 ;
        RECT  3.330 0.585 3.490 1.095 ;
        RECT  2.760 0.585 3.330 0.745 ;
        RECT  3.130 1.430 3.290 2.590 ;
        RECT  2.950 2.950 3.280 3.110 ;
        RECT  3.100 1.430 3.130 1.590 ;
        RECT  2.940 0.935 3.100 1.590 ;
        RECT  2.790 1.940 2.950 3.110 ;
        RECT  2.760 1.940 2.790 2.100 ;
        RECT  2.600 0.585 2.760 2.100 ;
        RECT  2.450 2.420 2.610 3.105 ;
        RECT  2.500 1.375 2.600 1.635 ;
        RECT  0.965 2.945 2.450 3.105 ;
        RECT  2.260 0.615 2.420 1.195 ;
        RECT  0.800 0.615 2.260 0.775 ;
        RECT  1.530 1.135 1.790 1.425 ;
        RECT  0.955 1.135 1.530 1.295 ;
        RECT  0.855 2.265 1.185 2.425 ;
        RECT  0.705 2.945 0.965 3.205 ;
        RECT  0.855 1.035 0.955 1.295 ;
        RECT  0.695 1.035 0.855 2.425 ;
        RECT  0.590 0.505 0.800 0.775 ;
        RECT  0.555 1.955 0.695 2.215 ;
        RECT  0.540 0.505 0.590 0.665 ;
    END
END SDFFXL

MACRO EDFFTRX4
    CLASS CORE ;
    FOREIGN EDFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.800 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 0.470 2.175 0.760 ;
        RECT  1.745 0.600 1.965 0.760 ;
        RECT  1.585 0.600 1.745 1.115 ;
        RECT  1.485 0.955 1.585 1.115 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.165 0.635 13.215 2.585 ;
        RECT  13.005 0.635 13.165 2.895 ;
        RECT  12.905 0.635 13.005 1.235 ;
        RECT  12.905 1.935 13.005 2.895 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.145 1.290 12.295 1.990 ;
        RECT  11.885 0.695 12.145 2.215 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 0.915 3.400 1.175 ;
        RECT  3.140 0.915 3.240 2.085 ;
        RECT  3.080 0.920 3.140 2.085 ;
        RECT  1.715 1.925 3.080 2.085 ;
        RECT  1.530 1.635 1.715 2.085 ;
        RECT  1.505 1.635 1.530 1.990 ;
        RECT  1.195 1.635 1.505 1.795 ;
        END
        ANTENNAGATEAREA     0.1729 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.290 4.015 1.605 ;
        RECT  3.420 1.355 3.805 1.605 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.190 0.335 1.875 ;
        END
        ANTENNAGATEAREA     0.2431 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.675 -0.250 13.800 0.250 ;
        RECT  13.415 -0.250 13.675 1.095 ;
        RECT  12.655 -0.250 13.415 0.250 ;
        RECT  12.395 -0.250 12.655 1.095 ;
        RECT  11.585 -0.250 12.395 0.250 ;
        RECT  11.585 0.495 11.635 0.755 ;
        RECT  11.425 -0.250 11.585 0.755 ;
        RECT  10.695 -0.250 11.425 0.250 ;
        RECT  11.375 0.495 11.425 0.755 ;
        RECT  10.435 -0.250 10.695 0.405 ;
        RECT  9.075 -0.250 10.435 0.250 ;
        RECT  8.815 -0.250 9.075 0.925 ;
        RECT  7.190 -0.250 8.815 0.250 ;
        RECT  6.930 -0.250 7.190 0.950 ;
        RECT  5.475 -0.250 6.930 0.250 ;
        RECT  5.215 -0.250 5.475 0.900 ;
        RECT  1.275 -0.250 5.215 0.250 ;
        RECT  0.675 -0.250 1.275 0.405 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.675 3.440 13.800 3.940 ;
        RECT  13.415 2.255 13.675 3.940 ;
        RECT  12.655 3.440 13.415 3.940 ;
        RECT  12.395 2.810 12.655 3.940 ;
        RECT  11.635 3.440 12.395 3.940 ;
        RECT  11.375 2.810 11.635 3.940 ;
        RECT  10.545 3.440 11.375 3.940 ;
        RECT  10.285 2.215 10.545 3.940 ;
        RECT  8.705 3.440 10.285 3.940 ;
        RECT  8.445 3.040 8.705 3.940 ;
        RECT  6.870 3.440 8.445 3.940 ;
        RECT  6.610 3.285 6.870 3.940 ;
        RECT  5.210 3.440 6.610 3.940 ;
        RECT  4.950 3.285 5.210 3.940 ;
        RECT  2.775 3.440 4.950 3.940 ;
        RECT  2.515 3.285 2.775 3.940 ;
        RECT  0.895 3.440 2.515 3.940 ;
        RECT  0.635 2.955 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.725 1.415 12.825 1.675 ;
        RECT  12.565 1.415 12.725 2.555 ;
        RECT  11.705 2.395 12.565 2.555 ;
        RECT  11.545 1.055 11.705 2.555 ;
        RECT  10.975 1.055 11.545 1.215 ;
        RECT  11.125 2.095 11.545 2.255 ;
        RECT  11.100 1.415 11.360 1.675 ;
        RECT  10.865 1.860 11.125 2.905 ;
        RECT  10.795 1.415 11.100 1.575 ;
        RECT  10.450 1.860 10.865 2.020 ;
        RECT  10.635 0.995 10.795 1.575 ;
        RECT  9.895 0.995 10.635 1.155 ;
        RECT  10.290 1.585 10.450 2.020 ;
        RECT  10.190 1.585 10.290 1.980 ;
        RECT  10.070 1.820 10.190 1.980 ;
        RECT  9.415 0.430 10.155 0.590 ;
        RECT  9.910 1.820 10.070 2.875 ;
        RECT  9.225 2.715 9.910 2.875 ;
        RECT  9.845 0.895 9.895 1.155 ;
        RECT  9.725 0.895 9.845 1.640 ;
        RECT  9.665 0.895 9.725 2.365 ;
        RECT  9.635 0.895 9.665 2.535 ;
        RECT  9.565 1.480 9.635 2.535 ;
        RECT  8.075 1.480 9.565 1.640 ;
        RECT  9.405 2.205 9.565 2.535 ;
        RECT  9.255 0.430 9.415 1.300 ;
        RECT  7.855 2.205 9.405 2.365 ;
        RECT  9.125 1.820 9.385 2.020 ;
        RECT  8.635 1.140 9.255 1.300 ;
        RECT  9.065 2.700 9.225 2.875 ;
        RECT  7.780 1.860 9.125 2.020 ;
        RECT  8.265 2.700 9.065 2.860 ;
        RECT  8.475 0.470 8.635 1.300 ;
        RECT  7.685 0.470 8.475 0.630 ;
        RECT  8.105 2.700 8.265 3.105 ;
        RECT  8.075 0.810 8.135 0.970 ;
        RECT  6.400 2.945 8.105 3.105 ;
        RECT  7.915 0.810 8.075 1.640 ;
        RECT  7.875 0.810 7.915 0.970 ;
        RECT  7.595 2.205 7.855 2.620 ;
        RECT  7.685 1.765 7.780 2.025 ;
        RECT  7.525 0.470 7.685 2.025 ;
        RECT  7.520 1.765 7.525 2.025 ;
        RECT  6.845 1.865 7.520 2.025 ;
        RECT  6.685 1.185 6.845 2.760 ;
        RECT  6.060 2.600 6.685 2.760 ;
        RECT  6.505 0.840 6.680 1.000 ;
        RECT  6.345 0.430 6.505 2.420 ;
        RECT  6.240 2.945 6.400 3.220 ;
        RECT  6.160 0.430 6.345 0.590 ;
        RECT  6.060 2.260 6.345 2.420 ;
        RECT  5.615 3.060 6.240 3.220 ;
        RECT  5.870 1.490 6.130 1.750 ;
        RECT  5.800 2.600 6.060 2.880 ;
        RECT  5.870 0.970 5.990 1.255 ;
        RECT  5.830 0.970 5.870 2.420 ;
        RECT  5.710 1.090 5.830 2.420 ;
        RECT  4.290 2.600 5.800 2.760 ;
        RECT  5.270 1.090 5.710 1.255 ;
        RECT  5.520 2.260 5.710 2.420 ;
        RECT  5.455 2.940 5.615 3.220 ;
        RECT  5.320 1.815 5.480 2.075 ;
        RECT  4.630 2.940 5.455 3.100 ;
        RECT  4.715 1.915 5.320 2.075 ;
        RECT  5.010 1.090 5.270 1.595 ;
        RECT  4.590 0.860 4.715 2.310 ;
        RECT  4.470 2.940 4.630 3.220 ;
        RECT  4.555 0.810 4.590 2.310 ;
        RECT  4.330 0.810 4.555 1.070 ;
        RECT  4.235 2.150 4.555 2.310 ;
        RECT  3.115 3.060 4.470 3.220 ;
        RECT  4.215 1.310 4.375 1.970 ;
        RECT  3.895 2.600 4.290 2.880 ;
        RECT  4.075 2.150 4.235 2.415 ;
        RECT  3.895 1.810 4.215 1.970 ;
        RECT  3.790 0.545 4.050 0.805 ;
        RECT  3.735 1.810 3.895 2.880 ;
        RECT  2.900 0.575 3.790 0.735 ;
        RECT  3.650 2.265 3.735 2.880 ;
        RECT  1.655 2.265 3.650 2.425 ;
        RECT  3.310 2.605 3.470 2.865 ;
        RECT  1.995 2.605 3.310 2.765 ;
        RECT  2.955 2.945 3.115 3.220 ;
        RECT  2.335 2.945 2.955 3.105 ;
        RECT  2.740 0.575 2.900 1.100 ;
        RECT  2.740 1.295 2.900 1.655 ;
        RECT  2.035 0.940 2.740 1.100 ;
        RECT  1.305 1.295 2.740 1.455 ;
        RECT  2.175 2.945 2.335 3.260 ;
        RECT  1.820 3.100 2.175 3.260 ;
        RECT  1.835 2.605 1.995 2.920 ;
        RECT  1.405 2.760 1.835 2.920 ;
        RECT  1.495 2.265 1.655 2.575 ;
        RECT  0.675 2.415 1.495 2.575 ;
        RECT  1.145 2.760 1.405 3.065 ;
        RECT  1.155 1.975 1.315 2.235 ;
        RECT  1.145 1.035 1.305 1.455 ;
        RECT  1.015 1.975 1.155 2.135 ;
        RECT  1.015 1.085 1.145 1.455 ;
        RECT  0.855 1.085 1.015 2.135 ;
        RECT  0.515 0.850 0.675 2.575 ;
        RECT  0.385 0.850 0.515 1.010 ;
        RECT  0.385 2.125 0.515 2.575 ;
        RECT  0.125 0.750 0.385 1.010 ;
        RECT  0.125 2.125 0.385 3.065 ;
    END
END EDFFTRX4

MACRO EDFFTRX2
    CLASS CORE ;
    FOREIGN EDFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 0.695 1.715 1.095 ;
        RECT  1.255 0.695 1.555 0.855 ;
        RECT  1.045 0.470 1.255 0.855 ;
        END
        ANTENNAGATEAREA     0.0611 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.710 0.695 11.835 2.585 ;
        RECT  11.550 0.695 11.710 3.025 ;
        RECT  11.435 2.085 11.550 3.025 ;
        END
        ANTENNADIFFAREA     0.7442 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.720 2.110 10.915 2.400 ;
        RECT  10.600 0.495 10.720 2.400 ;
        RECT  10.560 0.495 10.600 2.765 ;
        RECT  10.460 0.495 10.560 0.755 ;
        RECT  10.340 2.165 10.560 2.765 ;
        END
        ANTENNADIFFAREA     0.6614 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.105 1.095 3.350 1.355 ;
        RECT  2.945 1.095 3.105 1.860 ;
        RECT  2.560 1.700 2.945 1.860 ;
        RECT  2.300 1.635 2.560 1.895 ;
        RECT  2.150 1.700 2.300 1.895 ;
        RECT  1.715 1.700 2.150 1.860 ;
        RECT  1.505 1.635 1.715 1.990 ;
        RECT  1.195 1.635 1.505 1.795 ;
        END
        ANTENNAGATEAREA     0.1196 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.285 1.555 3.555 2.085 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.190 0.335 1.875 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.260 -0.250 11.960 0.250 ;
        RECT  11.000 -0.250 11.260 1.140 ;
        RECT  9.770 -0.250 11.000 0.250 ;
        RECT  9.510 -0.250 9.770 0.405 ;
        RECT  8.550 -0.250 9.510 0.250 ;
        RECT  8.290 -0.250 8.550 0.575 ;
        RECT  6.790 -0.250 8.290 0.250 ;
        RECT  6.530 -0.250 6.790 0.655 ;
        RECT  5.435 -0.250 6.530 0.250 ;
        RECT  5.275 -0.250 5.435 0.700 ;
        RECT  0.850 -0.250 5.275 0.250 ;
        RECT  0.590 -0.250 0.850 0.405 ;
        RECT  0.000 -0.250 0.590 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.140 3.440 11.960 3.940 ;
        RECT  10.880 3.285 11.140 3.940 ;
        RECT  9.540 3.440 10.880 3.940 ;
        RECT  9.280 3.285 9.540 3.940 ;
        RECT  8.430 3.440 9.280 3.940 ;
        RECT  8.170 3.285 8.430 3.940 ;
        RECT  6.720 3.440 8.170 3.940 ;
        RECT  6.460 3.285 6.720 3.940 ;
        RECT  5.155 3.440 6.460 3.940 ;
        RECT  4.895 3.285 5.155 3.940 ;
        RECT  2.775 3.440 4.895 3.940 ;
        RECT  2.515 3.285 2.775 3.940 ;
        RECT  0.935 3.440 2.515 3.940 ;
        RECT  0.675 2.895 0.935 3.940 ;
        RECT  0.000 3.440 0.675 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.255 1.560 11.370 1.820 ;
        RECT  11.095 1.560 11.255 3.105 ;
        RECT  10.090 2.945 11.095 3.105 ;
        RECT  10.200 1.015 10.360 1.980 ;
        RECT  10.060 1.015 10.200 1.275 ;
        RECT  10.090 1.820 10.200 1.980 ;
        RECT  9.930 1.820 10.090 3.105 ;
        RECT  9.030 1.470 10.020 1.630 ;
        RECT  9.830 1.965 9.930 2.625 ;
        RECT  9.245 1.965 9.830 2.125 ;
        RECT  9.145 1.810 9.245 2.125 ;
        RECT  9.130 0.435 9.230 0.695 ;
        RECT  8.985 1.810 9.145 3.105 ;
        RECT  8.970 0.435 9.130 0.915 ;
        RECT  8.800 1.095 9.030 1.630 ;
        RECT  6.280 2.945 8.985 3.105 ;
        RECT  8.045 0.755 8.970 0.915 ;
        RECT  8.770 1.095 8.800 2.765 ;
        RECT  8.640 1.425 8.770 2.765 ;
        RECT  7.670 1.425 8.640 1.585 ;
        RECT  8.540 2.360 8.640 2.765 ;
        RECT  7.580 2.360 8.540 2.520 ;
        RECT  7.885 0.545 8.045 0.915 ;
        RECT  7.230 0.545 7.885 0.705 ;
        RECT  7.510 0.885 7.670 1.585 ;
        RECT  7.320 2.360 7.580 2.765 ;
        RECT  7.410 0.885 7.510 1.145 ;
        RECT  7.230 1.915 7.410 2.175 ;
        RECT  7.070 0.545 7.230 2.175 ;
        RECT  6.580 2.015 7.070 2.175 ;
        RECT  6.420 1.305 6.580 2.760 ;
        RECT  6.390 1.305 6.420 1.570 ;
        RECT  5.935 2.600 6.420 2.760 ;
        RECT  6.120 2.945 6.280 3.260 ;
        RECT  6.210 0.555 6.245 0.815 ;
        RECT  6.210 2.160 6.240 2.420 ;
        RECT  6.050 0.430 6.210 2.420 ;
        RECT  5.495 3.100 6.120 3.260 ;
        RECT  5.985 0.430 6.050 0.815 ;
        RECT  5.615 0.430 5.985 0.590 ;
        RECT  5.675 2.600 5.935 2.920 ;
        RECT  5.710 1.090 5.870 2.420 ;
        RECT  5.680 1.090 5.710 1.350 ;
        RECT  5.645 1.790 5.710 2.420 ;
        RECT  4.930 1.090 5.680 1.255 ;
        RECT  4.315 2.600 5.675 2.760 ;
        RECT  5.570 2.160 5.645 2.420 ;
        RECT  5.335 2.940 5.495 3.260 ;
        RECT  5.200 1.960 5.360 2.250 ;
        RECT  4.655 2.940 5.335 3.100 ;
        RECT  4.430 2.090 5.200 2.250 ;
        RECT  4.770 1.090 4.930 1.910 ;
        RECT  4.670 1.650 4.770 1.910 ;
        RECT  4.495 2.940 4.655 3.220 ;
        RECT  4.430 0.645 4.600 0.905 ;
        RECT  3.245 3.060 4.495 3.220 ;
        RECT  4.340 0.645 4.430 2.310 ;
        RECT  4.270 0.650 4.340 2.310 ;
        RECT  4.055 2.600 4.315 2.870 ;
        RECT  4.265 2.150 4.270 2.310 ;
        RECT  4.105 2.150 4.265 2.415 ;
        RECT  3.930 1.090 4.090 1.970 ;
        RECT  3.925 2.600 4.055 2.760 ;
        RECT  3.770 0.645 4.030 0.905 ;
        RECT  3.925 1.810 3.930 1.970 ;
        RECT  3.765 1.810 3.925 2.760 ;
        RECT  2.085 0.745 3.770 0.905 ;
        RECT  1.655 2.265 3.765 2.425 ;
        RECT  3.425 2.605 3.585 2.865 ;
        RECT  1.995 2.605 3.425 2.765 ;
        RECT  3.085 2.945 3.245 3.220 ;
        RECT  2.335 2.945 3.085 3.105 ;
        RECT  2.605 1.150 2.765 1.455 ;
        RECT  1.345 1.295 2.605 1.455 ;
        RECT  2.175 2.945 2.335 3.260 ;
        RECT  1.945 3.100 2.175 3.260 ;
        RECT  1.925 0.745 2.085 1.115 ;
        RECT  1.835 2.605 1.995 2.915 ;
        RECT  1.525 2.755 1.835 2.915 ;
        RECT  1.495 2.265 1.655 2.575 ;
        RECT  1.265 2.755 1.525 3.045 ;
        RECT  0.675 2.415 1.495 2.575 ;
        RECT  1.185 1.035 1.345 1.455 ;
        RECT  1.155 1.975 1.315 2.235 ;
        RECT  1.015 1.085 1.185 1.455 ;
        RECT  1.015 1.975 1.155 2.135 ;
        RECT  0.855 1.085 1.015 2.135 ;
        RECT  0.515 0.850 0.675 2.575 ;
        RECT  0.385 0.850 0.515 1.010 ;
        RECT  0.125 2.055 0.515 2.315 ;
        RECT  0.125 0.750 0.385 1.010 ;
    END
END EDFFTRX2

MACRO EDFFTRX1
    CLASS CORE ;
    FOREIGN EDFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.685 0.855 1.715 1.115 ;
        RECT  1.525 0.695 1.685 1.115 ;
        RECT  1.255 0.695 1.525 0.855 ;
        RECT  1.045 0.470 1.255 0.855 ;
        END
        ANTENNAGATEAREA     0.0390 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.975 1.105 9.995 2.595 ;
        RECT  9.765 1.035 9.975 2.595 ;
        RECT  9.715 1.035 9.765 1.295 ;
        RECT  9.715 1.995 9.765 2.595 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.375 0.665 9.535 2.810 ;
        RECT  9.325 0.665 9.375 0.945 ;
        RECT  9.325 2.335 9.375 2.810 ;
        RECT  8.960 0.665 9.325 0.825 ;
        RECT  9.075 2.595 9.325 2.755 ;
        RECT  9.065 2.595 9.075 2.995 ;
        RECT  8.805 2.595 9.065 3.195 ;
        RECT  8.700 0.565 8.960 0.825 ;
        END
        ANTENNADIFFAREA     0.3626 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.105 1.095 3.350 1.355 ;
        RECT  2.945 1.095 3.105 1.860 ;
        RECT  2.560 1.700 2.945 1.860 ;
        RECT  2.150 1.700 2.560 1.960 ;
        RECT  1.715 1.800 2.150 1.960 ;
        RECT  1.505 1.635 1.715 1.990 ;
        RECT  1.195 1.635 1.505 1.795 ;
        END
        ANTENNAGATEAREA     0.0936 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.285 1.555 3.555 2.085 ;
        END
        ANTENNAGATEAREA     0.0442 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.190 0.335 1.875 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.500 -0.250 10.120 0.250 ;
        RECT  9.240 -0.250 9.500 0.405 ;
        RECT  8.410 -0.250 9.240 0.250 ;
        RECT  8.150 -0.250 8.410 0.405 ;
        RECT  6.790 -0.250 8.150 0.250 ;
        RECT  6.530 -0.250 6.790 0.800 ;
        RECT  5.435 -0.250 6.530 0.250 ;
        RECT  5.275 -0.250 5.435 0.700 ;
        RECT  0.850 -0.250 5.275 0.250 ;
        RECT  0.590 -0.250 0.850 0.405 ;
        RECT  0.000 -0.250 0.590 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.575 3.440 10.120 3.940 ;
        RECT  9.315 3.285 9.575 3.940 ;
        RECT  8.525 3.440 9.315 3.940 ;
        RECT  8.265 2.935 8.525 3.940 ;
        RECT  8.195 3.285 8.265 3.940 ;
        RECT  6.720 3.440 8.195 3.940 ;
        RECT  6.460 3.285 6.720 3.940 ;
        RECT  5.155 3.440 6.460 3.940 ;
        RECT  4.895 3.285 5.155 3.940 ;
        RECT  2.775 3.440 4.895 3.940 ;
        RECT  2.515 3.285 2.775 3.940 ;
        RECT  0.785 3.440 2.515 3.940 ;
        RECT  0.525 2.895 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.000 1.585 9.150 1.845 ;
        RECT  9.000 2.085 9.035 2.385 ;
        RECT  8.840 1.075 9.000 2.385 ;
        RECT  8.730 1.075 8.840 1.335 ;
        RECT  8.775 2.085 8.840 2.385 ;
        RECT  8.260 2.225 8.775 2.385 ;
        RECT  8.400 1.585 8.660 1.845 ;
        RECT  7.810 1.585 8.400 1.745 ;
        RECT  8.160 2.125 8.260 2.385 ;
        RECT  8.000 2.125 8.160 2.755 ;
        RECT  7.920 2.595 8.000 2.755 ;
        RECT  7.760 2.595 7.920 3.105 ;
        RECT  7.150 0.430 7.810 0.590 ;
        RECT  7.650 0.970 7.810 2.415 ;
        RECT  6.280 2.945 7.760 3.105 ;
        RECT  7.410 0.970 7.650 1.230 ;
        RECT  7.580 2.255 7.650 2.415 ;
        RECT  7.420 2.255 7.580 2.705 ;
        RECT  7.150 1.815 7.470 2.075 ;
        RECT  7.320 2.445 7.420 2.705 ;
        RECT  6.990 0.430 7.150 2.075 ;
        RECT  6.580 1.915 6.990 2.075 ;
        RECT  6.420 1.340 6.580 2.760 ;
        RECT  6.390 1.340 6.420 1.600 ;
        RECT  5.935 2.600 6.420 2.760 ;
        RECT  6.120 2.945 6.280 3.260 ;
        RECT  6.210 2.160 6.240 2.420 ;
        RECT  6.050 0.430 6.210 2.420 ;
        RECT  5.495 3.100 6.120 3.260 ;
        RECT  6.035 0.430 6.050 0.780 ;
        RECT  5.615 0.430 6.035 0.590 ;
        RECT  5.675 2.600 5.935 2.920 ;
        RECT  5.710 1.030 5.870 2.420 ;
        RECT  4.930 1.090 5.710 1.255 ;
        RECT  5.695 1.650 5.710 1.910 ;
        RECT  5.570 2.160 5.710 2.420 ;
        RECT  4.315 2.600 5.675 2.760 ;
        RECT  5.335 2.940 5.495 3.260 ;
        RECT  5.200 1.960 5.360 2.250 ;
        RECT  4.655 2.940 5.335 3.100 ;
        RECT  4.430 2.090 5.200 2.250 ;
        RECT  4.770 1.090 4.930 1.910 ;
        RECT  4.670 1.650 4.770 1.910 ;
        RECT  4.495 2.940 4.655 3.220 ;
        RECT  4.430 0.650 4.600 0.910 ;
        RECT  3.245 3.060 4.495 3.220 ;
        RECT  4.270 0.650 4.430 2.310 ;
        RECT  3.925 2.600 4.315 2.870 ;
        RECT  4.265 2.150 4.270 2.310 ;
        RECT  4.105 2.150 4.265 2.415 ;
        RECT  3.930 1.090 4.090 1.970 ;
        RECT  3.770 0.650 4.030 0.910 ;
        RECT  3.925 1.810 3.930 1.970 ;
        RECT  3.765 1.810 3.925 2.870 ;
        RECT  2.085 0.750 3.770 0.910 ;
        RECT  1.655 2.265 3.765 2.425 ;
        RECT  3.425 2.605 3.585 2.865 ;
        RECT  1.995 2.605 3.425 2.765 ;
        RECT  3.085 2.945 3.245 3.220 ;
        RECT  2.335 2.945 3.085 3.105 ;
        RECT  2.605 1.220 2.765 1.480 ;
        RECT  1.345 1.295 2.605 1.455 ;
        RECT  2.175 2.945 2.335 3.260 ;
        RECT  1.945 3.100 2.175 3.260 ;
        RECT  1.925 0.750 2.085 1.110 ;
        RECT  1.835 2.605 1.995 2.915 ;
        RECT  1.365 2.755 1.835 2.915 ;
        RECT  1.495 2.265 1.655 2.575 ;
        RECT  0.675 2.415 1.495 2.575 ;
        RECT  1.105 2.755 1.365 3.045 ;
        RECT  1.185 1.035 1.345 1.455 ;
        RECT  1.155 1.975 1.315 2.235 ;
        RECT  1.015 1.085 1.185 1.455 ;
        RECT  1.015 1.975 1.155 2.135 ;
        RECT  0.855 1.085 1.015 2.135 ;
        RECT  0.515 0.850 0.675 2.575 ;
        RECT  0.385 0.850 0.515 1.010 ;
        RECT  0.125 2.055 0.515 2.315 ;
        RECT  0.125 0.750 0.385 1.010 ;
    END
END EDFFTRX1

MACRO EDFFTRXL
    CLASS CORE ;
    FOREIGN EDFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.685 0.855 1.715 1.115 ;
        RECT  1.525 0.695 1.685 1.115 ;
        RECT  1.255 0.695 1.525 0.855 ;
        RECT  1.045 0.470 1.255 0.855 ;
        END
        ANTENNAGATEAREA     0.0741 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.945 1.290 9.995 2.215 ;
        RECT  9.785 1.035 9.945 2.215 ;
        RECT  9.735 1.955 9.785 2.215 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.485 0.625 9.535 2.400 ;
        RECT  9.375 0.625 9.485 2.630 ;
        RECT  9.325 0.625 9.375 0.945 ;
        RECT  9.325 2.110 9.375 2.630 ;
        RECT  8.990 0.625 9.325 0.785 ;
        RECT  9.065 2.470 9.325 2.630 ;
        RECT  8.805 2.470 9.065 2.730 ;
        RECT  8.730 0.525 8.990 0.785 ;
        END
        ANTENNADIFFAREA     0.2312 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.105 1.120 3.350 1.380 ;
        RECT  2.945 1.120 3.105 1.815 ;
        RECT  2.560 1.655 2.945 1.815 ;
        RECT  2.175 1.655 2.560 1.915 ;
        RECT  1.965 1.635 2.175 1.990 ;
        RECT  1.195 1.635 1.965 1.795 ;
        END
        ANTENNAGATEAREA     0.1352 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.285 1.560 3.555 2.085 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.190 0.335 1.780 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.500 -0.250 10.120 0.250 ;
        RECT  9.240 -0.250 9.500 0.405 ;
        RECT  8.410 -0.250 9.240 0.250 ;
        RECT  8.150 -0.250 8.410 0.405 ;
        RECT  6.790 -0.250 8.150 0.250 ;
        RECT  6.530 -0.250 6.790 0.795 ;
        RECT  5.435 -0.250 6.530 0.250 ;
        RECT  5.275 -0.250 5.435 0.700 ;
        RECT  0.850 -0.250 5.275 0.250 ;
        RECT  0.590 -0.250 0.850 0.405 ;
        RECT  0.000 -0.250 0.590 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.575 3.440 10.120 3.940 ;
        RECT  9.315 2.895 9.575 3.940 ;
        RECT  8.490 3.440 9.315 3.940 ;
        RECT  8.230 2.895 8.490 3.940 ;
        RECT  6.720 3.440 8.230 3.940 ;
        RECT  6.460 3.285 6.720 3.940 ;
        RECT  5.155 3.440 6.460 3.940 ;
        RECT  4.895 3.285 5.155 3.940 ;
        RECT  2.805 3.440 4.895 3.940 ;
        RECT  2.545 3.285 2.805 3.940 ;
        RECT  0.815 3.440 2.545 3.940 ;
        RECT  0.555 2.895 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.000 1.405 9.150 1.665 ;
        RECT  9.000 1.955 9.065 2.215 ;
        RECT  8.840 1.035 9.000 2.215 ;
        RECT  8.730 1.035 8.840 1.295 ;
        RECT  8.805 1.955 8.840 2.215 ;
        RECT  8.260 2.055 8.805 2.215 ;
        RECT  8.400 1.475 8.660 1.735 ;
        RECT  7.810 1.525 8.400 1.685 ;
        RECT  8.160 1.955 8.260 2.215 ;
        RECT  8.000 1.955 8.160 2.715 ;
        RECT  7.920 2.555 8.000 2.715 ;
        RECT  7.760 2.555 7.920 3.105 ;
        RECT  7.150 0.430 7.810 0.590 ;
        RECT  7.650 0.965 7.810 2.375 ;
        RECT  6.280 2.945 7.760 3.105 ;
        RECT  7.410 0.965 7.650 1.225 ;
        RECT  7.580 2.215 7.650 2.375 ;
        RECT  7.420 2.215 7.580 2.600 ;
        RECT  7.150 1.865 7.470 2.025 ;
        RECT  7.320 2.340 7.420 2.600 ;
        RECT  6.990 0.430 7.150 2.025 ;
        RECT  6.680 1.865 6.990 2.025 ;
        RECT  6.520 1.340 6.680 2.760 ;
        RECT  6.420 1.340 6.520 1.600 ;
        RECT  5.935 2.600 6.520 2.760 ;
        RECT  6.210 2.160 6.290 2.420 ;
        RECT  6.120 2.945 6.280 3.260 ;
        RECT  6.210 0.430 6.245 0.780 ;
        RECT  6.050 0.430 6.210 2.420 ;
        RECT  5.495 3.100 6.120 3.260 ;
        RECT  5.985 0.430 6.050 0.780 ;
        RECT  6.030 2.160 6.050 2.420 ;
        RECT  5.615 0.430 5.985 0.590 ;
        RECT  5.675 2.600 5.935 2.920 ;
        RECT  5.825 1.035 5.870 1.295 ;
        RECT  5.825 1.650 5.855 1.980 ;
        RECT  5.710 1.035 5.825 2.420 ;
        RECT  5.665 1.090 5.710 2.420 ;
        RECT  4.315 2.600 5.675 2.760 ;
        RECT  4.945 1.090 5.665 1.255 ;
        RECT  5.570 2.160 5.665 2.420 ;
        RECT  5.335 2.940 5.495 3.260 ;
        RECT  5.200 1.960 5.360 2.420 ;
        RECT  4.655 2.940 5.335 3.100 ;
        RECT  4.430 2.260 5.200 2.420 ;
        RECT  4.785 1.090 4.945 1.910 ;
        RECT  4.720 1.640 4.785 1.910 ;
        RECT  4.670 1.640 4.720 1.900 ;
        RECT  4.495 2.940 4.655 3.220 ;
        RECT  4.430 0.670 4.600 0.930 ;
        RECT  3.245 3.060 4.495 3.220 ;
        RECT  4.270 0.670 4.430 2.420 ;
        RECT  3.925 2.600 4.315 2.870 ;
        RECT  4.105 2.150 4.270 2.420 ;
        RECT  3.930 1.090 4.090 1.970 ;
        RECT  3.770 0.640 4.030 0.910 ;
        RECT  3.925 1.810 3.930 1.970 ;
        RECT  3.765 1.810 3.925 2.870 ;
        RECT  2.085 0.750 3.770 0.910 ;
        RECT  1.685 2.265 3.765 2.425 ;
        RECT  3.425 2.605 3.585 2.865 ;
        RECT  2.025 2.605 3.425 2.765 ;
        RECT  3.085 2.945 3.245 3.220 ;
        RECT  2.365 2.945 3.085 3.105 ;
        RECT  2.605 1.175 2.765 1.455 ;
        RECT  1.345 1.295 2.605 1.455 ;
        RECT  2.205 2.945 2.365 3.260 ;
        RECT  1.945 3.100 2.205 3.260 ;
        RECT  1.925 0.750 2.085 1.065 ;
        RECT  1.865 2.605 2.025 2.915 ;
        RECT  1.365 2.755 1.865 2.915 ;
        RECT  1.525 2.265 1.685 2.575 ;
        RECT  0.675 2.415 1.525 2.575 ;
        RECT  1.105 2.755 1.365 3.065 ;
        RECT  1.185 1.035 1.345 1.455 ;
        RECT  1.185 1.975 1.345 2.235 ;
        RECT  1.015 1.085 1.185 1.455 ;
        RECT  1.015 1.975 1.185 2.135 ;
        RECT  0.855 1.085 1.015 2.135 ;
        RECT  0.515 0.850 0.675 2.575 ;
        RECT  0.385 0.850 0.515 1.010 ;
        RECT  0.125 1.975 0.515 2.235 ;
        RECT  0.125 0.750 0.385 1.010 ;
    END
END EDFFTRXL

MACRO EDFFX4
    CLASS CORE ;
    FOREIGN EDFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 1.515 13.675 2.595 ;
        RECT  13.615 0.900 13.660 2.595 ;
        RECT  13.600 0.900 13.615 3.030 ;
        RECT  13.420 0.590 13.600 3.030 ;
        RECT  13.340 0.590 13.420 1.190 ;
        RECT  13.355 2.090 13.420 3.030 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.535 1.890 12.595 2.405 ;
        RECT  12.535 0.590 12.580 1.190 ;
        RECT  12.375 0.590 12.535 2.405 ;
        RECT  12.320 0.590 12.375 1.190 ;
        RECT  12.335 1.700 12.375 2.405 ;
        RECT  12.085 1.700 12.335 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 2.715 0.830 3.050 ;
        RECT  0.585 2.715 0.795 3.220 ;
        RECT  0.570 2.715 0.585 3.050 ;
        END
        ANTENNAGATEAREA     0.1703 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.700 1.635 1.990 ;
        END
        ANTENNAGATEAREA     0.1209 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 1.675 5.170 1.935 ;
        RECT  4.725 1.675 4.935 1.990 ;
        RECT  4.715 1.675 4.725 1.885 ;
        END
        ANTENNAGATEAREA     0.2327 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.110 -0.250 14.260 0.250 ;
        RECT  13.850 -0.250 14.110 1.190 ;
        RECT  13.090 -0.250 13.850 0.250 ;
        RECT  12.830 -0.250 13.090 1.190 ;
        RECT  12.070 -0.250 12.830 0.250 ;
        RECT  11.810 -0.250 12.070 1.190 ;
        RECT  10.920 -0.250 11.810 0.250 ;
        RECT  10.660 -0.250 10.920 1.210 ;
        RECT  8.905 -0.250 10.660 0.250 ;
        RECT  8.645 -0.250 8.905 0.890 ;
        RECT  7.230 -0.250 8.645 0.250 ;
        RECT  6.970 -0.250 7.230 0.955 ;
        RECT  5.550 -0.250 6.970 0.250 ;
        RECT  5.290 -0.250 5.550 0.405 ;
        RECT  4.590 -0.250 5.290 0.250 ;
        RECT  4.330 -0.250 4.590 0.405 ;
        RECT  2.270 -0.250 4.330 0.250 ;
        RECT  2.010 -0.250 2.270 0.730 ;
        RECT  0.405 -0.250 2.010 0.250 ;
        RECT  0.145 -0.250 0.405 1.295 ;
        RECT  0.000 -0.250 0.145 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.125 3.440 14.260 3.940 ;
        RECT  13.865 2.210 14.125 3.940 ;
        RECT  13.105 3.440 13.865 3.940 ;
        RECT  12.845 2.930 13.105 3.940 ;
        RECT  12.085 3.440 12.845 3.940 ;
        RECT  11.825 2.935 12.085 3.940 ;
        RECT  11.035 3.440 11.825 3.940 ;
        RECT  10.775 2.550 11.035 3.940 ;
        RECT  9.060 3.440 10.775 3.940 ;
        RECT  8.800 3.285 9.060 3.940 ;
        RECT  7.335 3.440 8.800 3.940 ;
        RECT  7.075 3.285 7.335 3.940 ;
        RECT  5.675 3.440 7.075 3.940 ;
        RECT  5.415 3.285 5.675 3.940 ;
        RECT  4.610 3.440 5.415 3.940 ;
        RECT  4.350 3.285 4.610 3.940 ;
        RECT  2.265 3.440 4.350 3.940 ;
        RECT  2.005 2.735 2.265 3.940 ;
        RECT  0.390 3.440 2.005 3.940 ;
        RECT  0.130 2.190 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.085 1.505 13.195 1.810 ;
        RECT  13.035 1.505 13.085 2.745 ;
        RECT  12.925 1.650 13.035 2.745 ;
        RECT  11.575 2.585 12.925 2.745 ;
        RECT  11.415 2.085 11.575 3.025 ;
        RECT  11.415 0.575 11.430 1.175 ;
        RECT  11.315 0.575 11.415 3.025 ;
        RECT  11.255 0.575 11.315 2.335 ;
        RECT  11.170 0.575 11.255 1.175 ;
        RECT  10.600 2.175 11.255 2.335 ;
        RECT  10.790 1.550 11.050 1.940 ;
        RECT  10.480 1.745 10.790 1.940 ;
        RECT  10.595 2.130 10.600 2.390 ;
        RECT  10.440 2.130 10.595 3.105 ;
        RECT  10.320 0.715 10.480 1.940 ;
        RECT  10.435 2.180 10.440 3.105 ;
        RECT  4.135 2.945 10.435 3.105 ;
        RECT  9.780 0.715 10.320 0.875 ;
        RECT  10.255 1.780 10.320 1.940 ;
        RECT  10.095 1.780 10.255 2.540 ;
        RECT  9.980 1.065 10.140 1.595 ;
        RECT  9.960 2.380 10.095 2.540 ;
        RECT  9.915 1.435 9.980 1.595 ;
        RECT  9.700 2.380 9.960 2.755 ;
        RECT  9.755 1.435 9.915 2.075 ;
        RECT  9.730 0.715 9.780 1.110 ;
        RECT  8.370 1.915 9.755 2.075 ;
        RECT  9.520 0.715 9.730 1.230 ;
        RECT  8.150 2.380 9.700 2.540 ;
        RECT  9.300 1.410 9.570 1.590 ;
        RECT  8.050 1.070 9.520 1.230 ;
        RECT  7.880 1.410 9.300 1.570 ;
        RECT  8.110 1.750 8.370 2.075 ;
        RECT  7.990 2.330 8.150 2.590 ;
        RECT  7.810 1.915 8.110 2.075 ;
        RECT  7.840 0.845 8.050 1.230 ;
        RECT  7.670 1.410 7.880 1.615 ;
        RECT  7.790 0.845 7.840 1.105 ;
        RECT  7.650 1.915 7.810 2.760 ;
        RECT  7.490 1.455 7.670 1.615 ;
        RECT  4.150 2.600 7.650 2.760 ;
        RECT  7.465 1.135 7.490 1.615 ;
        RECT  7.305 1.135 7.465 2.415 ;
        RECT  6.720 1.135 7.305 1.295 ;
        RECT  6.500 2.255 7.305 2.415 ;
        RECT  6.960 1.515 7.120 1.775 ;
        RECT  6.235 1.570 6.960 1.730 ;
        RECT  6.620 0.775 6.720 1.295 ;
        RECT  6.460 0.585 6.620 1.295 ;
        RECT  4.130 0.585 6.460 0.745 ;
        RECT  6.075 1.175 6.235 2.355 ;
        RECT  6.070 1.175 6.075 1.335 ;
        RECT  4.500 2.195 6.075 2.355 ;
        RECT  5.810 1.075 6.070 1.335 ;
        RECT  5.585 1.675 5.845 1.935 ;
        RECT  5.560 1.675 5.585 1.835 ;
        RECT  5.400 0.925 5.560 1.835 ;
        RECT  3.700 0.925 5.400 1.085 ;
        RECT  4.435 1.270 4.970 1.430 ;
        RECT  4.340 2.140 4.500 2.400 ;
        RECT  4.275 1.270 4.435 1.615 ;
        RECT  4.015 1.455 4.275 1.615 ;
        RECT  4.015 2.245 4.150 2.760 ;
        RECT  3.975 2.945 4.135 3.215 ;
        RECT  3.970 0.485 4.130 0.745 ;
        RECT  3.990 1.455 4.015 2.760 ;
        RECT  3.855 1.455 3.990 2.405 ;
        RECT  2.775 3.055 3.975 3.215 ;
        RECT  3.640 0.485 3.970 0.645 ;
        RECT  3.205 1.455 3.855 1.615 ;
        RECT  3.805 2.245 3.855 2.405 ;
        RECT  3.585 2.585 3.805 2.845 ;
        RECT  3.600 0.835 3.700 1.095 ;
        RECT  3.440 0.835 3.600 1.275 ;
        RECT  3.545 1.875 3.585 2.845 ;
        RECT  3.425 1.875 3.545 2.745 ;
        RECT  3.025 1.115 3.440 1.275 ;
        RECT  3.025 1.875 3.425 2.035 ;
        RECT  3.120 2.565 3.220 2.825 ;
        RECT  2.900 0.675 3.160 0.935 ;
        RECT  2.960 2.395 3.120 2.825 ;
        RECT  2.865 1.115 3.025 2.035 ;
        RECT  1.575 2.395 2.960 2.555 ;
        RECT  2.680 0.775 2.900 0.935 ;
        RECT  2.520 0.775 2.680 1.070 ;
        RECT  1.615 0.910 2.520 1.070 ;
        RECT  2.175 1.255 2.480 1.415 ;
        RECT  2.015 1.255 2.175 2.205 ;
        RECT  0.975 1.255 2.015 1.415 ;
        RECT  1.855 2.045 2.015 2.205 ;
        RECT  1.455 0.625 1.615 1.070 ;
        RECT  1.445 2.395 1.575 2.865 ;
        RECT  1.370 0.625 1.455 0.785 ;
        RECT  1.415 2.395 1.445 2.965 ;
        RECT  1.185 2.705 1.415 2.965 ;
        RECT  1.110 0.525 1.370 0.785 ;
        RECT  0.855 1.035 0.975 1.415 ;
        RECT  0.855 2.190 0.970 2.450 ;
        RECT  0.695 1.035 0.855 2.450 ;
    END
END EDFFX4

MACRO EDFFX2
    CLASS CORE ;
    FOREIGN EDFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.165 0.590 11.375 3.030 ;
        RECT  11.115 0.590 11.165 1.190 ;
        RECT  11.115 2.090 11.165 3.030 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.355 1.515 10.455 2.175 ;
        RECT  10.310 1.515 10.355 2.335 ;
        RECT  10.150 0.490 10.310 2.335 ;
        RECT  10.050 0.490 10.150 0.750 ;
        RECT  10.095 2.075 10.150 2.335 ;
        END
        ANTENNADIFFAREA     0.5803 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.350 1.615 0.385 1.875 ;
        RECT  0.335 1.525 0.350 1.875 ;
        RECT  0.125 1.290 0.335 1.875 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 1.650 1.170 1.905 ;
        RECT  0.780 1.650 0.945 1.990 ;
        RECT  0.585 1.700 0.780 1.990 ;
        END
        ANTENNAGATEAREA     0.0676 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.675 4.590 1.935 ;
        RECT  4.265 1.675 4.475 1.990 ;
        RECT  4.100 1.675 4.265 1.885 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.865 -0.250 11.500 0.250 ;
        RECT  10.605 -0.250 10.865 1.190 ;
        RECT  9.500 -0.250 10.605 0.250 ;
        RECT  9.240 -0.250 9.500 0.405 ;
        RECT  8.240 -0.250 9.240 0.250 ;
        RECT  7.980 -0.250 8.240 0.405 ;
        RECT  6.510 -0.250 7.980 0.250 ;
        RECT  6.510 0.860 6.560 1.120 ;
        RECT  6.250 -0.250 6.510 1.120 ;
        RECT  4.900 -0.250 6.250 0.250 ;
        RECT  3.960 -0.250 4.900 0.655 ;
        RECT  1.800 -0.250 3.960 0.250 ;
        RECT  1.540 -0.250 1.800 0.745 ;
        RECT  0.385 -0.250 1.540 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.865 3.440 11.500 3.940 ;
        RECT  10.605 2.930 10.865 3.940 ;
        RECT  9.520 3.440 10.605 3.940 ;
        RECT  9.260 3.285 9.520 3.940 ;
        RECT  8.680 3.440 9.260 3.940 ;
        RECT  8.080 3.285 8.680 3.940 ;
        RECT  6.620 3.440 8.080 3.940 ;
        RECT  5.680 3.285 6.620 3.940 ;
        RECT  4.890 3.440 5.680 3.940 ;
        RECT  3.800 3.285 4.890 3.940 ;
        RECT  1.745 3.440 3.800 3.940 ;
        RECT  1.485 2.865 1.745 3.940 ;
        RECT  0.385 3.440 1.485 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.935 1.505 10.955 1.765 ;
        RECT  10.775 1.505 10.935 2.745 ;
        RECT  9.920 2.585 10.775 2.745 ;
        RECT  9.910 2.585 9.920 2.870 ;
        RECT  9.750 1.000 9.910 2.870 ;
        RECT  9.650 1.000 9.750 1.260 ;
        RECT  9.660 2.530 9.750 2.870 ;
        RECT  9.115 2.530 9.660 2.690 ;
        RECT  9.205 1.550 9.570 1.810 ;
        RECT  9.045 1.100 9.205 2.310 ;
        RECT  8.955 2.530 9.115 3.125 ;
        RECT  8.610 1.100 9.045 1.260 ;
        RECT  8.780 2.150 9.045 2.310 ;
        RECT  8.855 2.865 8.955 3.125 ;
        RECT  3.460 2.890 8.855 3.050 ;
        RECT  8.695 1.480 8.795 1.740 ;
        RECT  8.680 2.150 8.780 2.410 ;
        RECT  8.535 1.480 8.695 1.940 ;
        RECT  8.520 2.150 8.680 2.625 ;
        RECT  8.350 1.000 8.610 1.260 ;
        RECT  7.650 1.780 8.535 1.940 ;
        RECT  7.430 2.465 8.520 2.625 ;
        RECT  7.380 1.025 8.350 1.185 ;
        RECT  7.485 1.780 7.650 2.190 ;
        RECT  7.330 1.410 7.550 1.570 ;
        RECT  7.090 1.930 7.485 2.190 ;
        RECT  7.270 2.415 7.430 2.675 ;
        RECT  7.170 0.795 7.380 1.185 ;
        RECT  6.950 1.400 7.330 1.570 ;
        RECT  7.120 0.795 7.170 1.055 ;
        RECT  7.050 1.930 7.090 2.705 ;
        RECT  6.930 2.030 7.050 2.705 ;
        RECT  6.745 1.400 6.950 1.560 ;
        RECT  4.420 2.545 6.930 2.705 ;
        RECT  6.585 1.330 6.745 2.360 ;
        RECT  5.930 1.330 6.585 1.560 ;
        RECT  6.150 2.200 6.585 2.360 ;
        RECT  6.240 1.745 6.400 2.005 ;
        RECT  5.565 1.795 6.240 1.955 ;
        RECT  5.885 2.170 6.150 2.360 ;
        RECT  5.770 0.565 5.930 1.560 ;
        RECT  5.480 0.565 5.770 0.725 ;
        RECT  5.405 1.225 5.565 2.330 ;
        RECT  5.220 0.465 5.480 0.725 ;
        RECT  5.210 1.225 5.405 1.385 ;
        RECT  3.800 2.170 5.405 2.330 ;
        RECT  5.055 1.675 5.215 1.935 ;
        RECT  4.950 1.675 5.055 1.835 ;
        RECT  4.790 0.880 4.950 1.835 ;
        RECT  3.260 0.880 4.790 1.040 ;
        RECT  4.160 2.510 4.420 2.705 ;
        RECT  3.745 1.225 4.270 1.385 ;
        RECT  3.460 2.545 4.160 2.705 ;
        RECT  3.640 1.810 3.800 2.330 ;
        RECT  3.585 1.225 3.745 1.605 ;
        RECT  3.320 1.445 3.585 1.605 ;
        RECT  3.320 2.245 3.460 2.705 ;
        RECT  3.300 2.890 3.460 3.215 ;
        RECT  3.300 1.445 3.320 2.705 ;
        RECT  3.160 1.445 3.300 2.455 ;
        RECT  2.170 3.055 3.300 3.215 ;
        RECT  3.160 0.750 3.260 1.040 ;
        RECT  3.000 0.750 3.160 1.265 ;
        RECT  2.720 1.445 3.160 1.605 ;
        RECT  2.940 2.655 3.105 2.815 ;
        RECT  2.540 1.105 3.000 1.265 ;
        RECT  2.780 1.875 2.940 2.815 ;
        RECT  2.540 1.875 2.780 2.035 ;
        RECT  2.155 0.765 2.690 0.925 ;
        RECT  2.385 2.525 2.545 2.850 ;
        RECT  2.380 1.105 2.540 2.035 ;
        RECT  1.200 2.525 2.385 2.685 ;
        RECT  1.995 0.765 2.155 1.085 ;
        RECT  1.640 1.265 2.010 1.525 ;
        RECT  1.245 0.925 1.995 1.085 ;
        RECT  1.480 1.265 1.640 2.345 ;
        RECT  0.825 1.265 1.480 1.425 ;
        RECT  1.285 2.085 1.480 2.345 ;
        RECT  0.555 2.185 1.285 2.345 ;
        RECT  1.085 0.570 1.245 1.085 ;
        RECT  1.040 2.525 1.200 2.805 ;
        RECT  0.640 0.570 1.085 0.730 ;
        RECT  0.895 2.645 1.040 2.805 ;
        RECT  0.635 2.645 0.895 2.905 ;
        RECT  0.665 1.030 0.825 1.425 ;
        RECT  0.565 1.030 0.665 1.290 ;
    END
END EDFFX2

MACRO EDFFX1
    CLASS CORE ;
    FOREIGN EDFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.485 1.105 9.535 2.825 ;
        RECT  9.325 0.975 9.485 2.825 ;
        RECT  9.275 2.225 9.325 2.825 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.075 0.675 9.145 2.075 ;
        RECT  8.985 0.675 9.075 2.815 ;
        RECT  8.865 0.675 8.985 0.945 ;
        RECT  8.915 1.915 8.985 2.815 ;
        RECT  8.865 2.330 8.915 2.815 ;
        RECT  8.595 0.675 8.865 0.835 ;
        RECT  8.615 2.655 8.865 2.815 ;
        RECT  8.580 2.655 8.615 2.995 ;
        RECT  8.335 0.575 8.595 0.835 ;
        RECT  8.370 2.655 8.580 3.070 ;
        RECT  8.320 2.810 8.370 3.070 ;
        END
        ANTENNADIFFAREA     0.3264 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.635 0.410 1.895 ;
        RECT  0.150 1.635 0.335 2.810 ;
        RECT  0.125 1.895 0.150 2.810 ;
        END
        ANTENNAGATEAREA     0.0923 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.665 2.415 1.925 ;
        RECT  2.015 1.290 2.175 1.925 ;
        RECT  1.965 1.290 2.015 1.580 ;
        END
        ANTENNAGATEAREA     0.0429 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.370 1.290 5.395 1.580 ;
        RECT  5.195 1.290 5.370 1.675 ;
        RECT  5.185 1.290 5.195 1.715 ;
        RECT  4.795 1.515 5.185 1.715 ;
        END
        ANTENNAGATEAREA     0.0832 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.135 -0.250 9.660 0.250 ;
        RECT  8.875 -0.250 9.135 0.405 ;
        RECT  8.045 -0.250 8.875 0.250 ;
        RECT  7.785 -0.250 8.045 0.405 ;
        RECT  6.455 -0.250 7.785 0.250 ;
        RECT  6.295 -0.250 6.455 0.625 ;
        RECT  5.095 -0.250 6.295 0.250 ;
        RECT  4.935 -0.250 5.095 0.690 ;
        RECT  4.065 -0.250 4.935 0.250 ;
        RECT  3.805 -0.250 4.065 0.895 ;
        RECT  1.865 -0.250 3.805 0.250 ;
        RECT  1.605 -0.250 1.865 0.405 ;
        RECT  0.385 -0.250 1.605 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.095 3.440 9.660 3.940 ;
        RECT  8.835 3.285 9.095 3.940 ;
        RECT  8.070 3.440 8.835 3.940 ;
        RECT  7.810 2.810 8.070 3.940 ;
        RECT  7.775 3.285 7.810 3.940 ;
        RECT  5.640 3.440 7.775 3.940 ;
        RECT  5.380 3.285 5.640 3.940 ;
        RECT  3.715 3.440 5.380 3.940 ;
        RECT  3.455 3.285 3.715 3.940 ;
        RECT  1.745 3.440 3.455 3.940 ;
        RECT  1.485 3.285 1.745 3.940 ;
        RECT  0.385 3.440 1.485 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.635 1.475 8.805 1.735 ;
        RECT  8.475 1.105 8.635 2.385 ;
        RECT  8.365 1.105 8.475 1.365 ;
        RECT  8.325 2.125 8.475 2.385 ;
        RECT  7.490 2.175 8.325 2.335 ;
        RECT  8.035 1.545 8.295 1.805 ;
        RECT  7.095 1.645 8.035 1.805 ;
        RECT  7.490 2.850 7.615 3.110 ;
        RECT  7.330 2.175 7.490 3.160 ;
        RECT  7.185 0.535 7.445 0.795 ;
        RECT  6.525 3.000 7.330 3.160 ;
        RECT  7.095 0.975 7.305 1.320 ;
        RECT  6.850 0.635 7.185 0.795 ;
        RECT  7.045 0.975 7.095 2.740 ;
        RECT  6.965 1.160 7.045 2.740 ;
        RECT  6.935 1.160 6.965 2.790 ;
        RECT  6.705 2.530 6.935 2.790 ;
        RECT  6.690 0.635 6.850 0.980 ;
        RECT  6.525 2.190 6.755 2.350 ;
        RECT  6.525 0.805 6.690 0.980 ;
        RECT  6.365 0.805 6.525 2.765 ;
        RECT  6.365 2.945 6.525 3.160 ;
        RECT  6.115 0.805 6.365 0.965 ;
        RECT  4.495 2.605 6.365 2.765 ;
        RECT  4.840 2.945 6.365 3.105 ;
        RECT  6.025 1.485 6.185 2.410 ;
        RECT  5.955 0.430 6.115 0.965 ;
        RECT  5.975 1.485 6.025 1.645 ;
        RECT  5.200 2.250 6.025 2.410 ;
        RECT  5.815 1.145 5.975 1.645 ;
        RECT  5.435 0.430 5.955 0.590 ;
        RECT  5.795 1.905 5.845 2.065 ;
        RECT  5.775 1.145 5.815 1.305 ;
        RECT  5.585 1.895 5.795 2.065 ;
        RECT  5.615 0.770 5.775 1.305 ;
        RECT  4.515 1.895 5.585 2.055 ;
        RECT  5.275 0.430 5.435 1.060 ;
        RECT  4.805 0.900 5.275 1.060 ;
        RECT  5.040 2.235 5.200 2.410 ;
        RECT  4.805 2.235 5.040 2.395 ;
        RECT  4.680 2.945 4.840 3.260 ;
        RECT  4.645 0.900 4.805 1.335 ;
        RECT  4.055 3.100 4.680 3.260 ;
        RECT  4.465 0.550 4.635 0.710 ;
        RECT  4.465 1.895 4.515 2.215 ;
        RECT  4.395 2.605 4.495 2.920 ;
        RECT  4.305 0.550 4.465 2.215 ;
        RECT  4.235 2.410 4.395 2.920 ;
        RECT  3.865 1.085 4.305 1.245 ;
        RECT  4.235 2.055 4.305 2.215 ;
        RECT  3.365 2.410 4.235 2.570 ;
        RECT  3.965 1.565 4.125 1.825 ;
        RECT  3.895 2.940 4.055 3.260 ;
        RECT  3.185 1.565 3.965 1.725 ;
        RECT  1.065 2.940 3.895 3.100 ;
        RECT  3.605 1.085 3.865 1.345 ;
        RECT  3.105 2.410 3.365 2.670 ;
        RECT  3.025 0.750 3.185 2.215 ;
        RECT  2.775 2.410 3.105 2.570 ;
        RECT  2.925 0.750 3.025 1.010 ;
        RECT  2.955 1.955 3.025 2.215 ;
        RECT  2.745 1.190 2.775 2.570 ;
        RECT  2.615 1.090 2.745 2.570 ;
        RECT  2.420 0.650 2.615 0.910 ;
        RECT  2.485 1.090 2.615 1.350 ;
        RECT  2.275 2.160 2.435 2.720 ;
        RECT  2.260 0.585 2.420 0.910 ;
        RECT  0.815 2.560 2.275 2.720 ;
        RECT  0.975 0.585 2.260 0.745 ;
        RECT  1.545 1.910 1.805 2.170 ;
        RECT  1.500 1.115 1.600 1.375 ;
        RECT  1.500 1.910 1.545 2.070 ;
        RECT  1.340 1.115 1.500 2.070 ;
        RECT  0.815 1.135 1.340 1.295 ;
        RECT  0.905 2.940 1.065 3.210 ;
        RECT  0.765 0.475 0.975 0.745 ;
        RECT  0.805 2.950 0.905 3.210 ;
        RECT  0.765 1.035 0.815 1.295 ;
        RECT  0.765 2.050 0.815 2.310 ;
        RECT  0.550 2.560 0.815 2.770 ;
        RECT  0.715 0.475 0.765 0.635 ;
        RECT  0.605 1.035 0.765 2.310 ;
        RECT  0.555 1.035 0.605 1.295 ;
        RECT  0.555 2.050 0.605 2.310 ;
    END
END EDFFX1

MACRO EDFFXL
    CLASS CORE ;
    FOREIGN EDFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.485 1.105 9.535 2.655 ;
        RECT  9.325 0.995 9.485 2.655 ;
        RECT  9.275 2.395 9.325 2.655 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.075 1.105 9.145 2.075 ;
        RECT  8.985 1.105 9.075 2.815 ;
        RECT  8.975 1.105 8.985 1.295 ;
        RECT  8.915 1.915 8.985 2.815 ;
        RECT  8.815 0.615 8.975 1.295 ;
        RECT  8.865 2.335 8.915 2.815 ;
        RECT  8.580 2.655 8.865 2.815 ;
        RECT  8.595 0.615 8.815 0.775 ;
        RECT  8.335 0.575 8.595 0.835 ;
        RECT  8.370 2.655 8.580 3.035 ;
        RECT  8.320 2.775 8.370 3.035 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.635 0.360 1.895 ;
        RECT  0.150 1.635 0.335 2.810 ;
        RECT  0.125 1.895 0.150 2.810 ;
        END
        ANTENNAGATEAREA     0.1313 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.195 1.960 2.335 2.120 ;
        RECT  2.175 1.355 2.195 2.120 ;
        RECT  2.035 1.290 2.175 2.120 ;
        RECT  1.965 1.290 2.035 1.580 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.370 1.290 5.395 1.580 ;
        RECT  5.195 1.290 5.370 1.675 ;
        RECT  5.185 1.290 5.195 1.715 ;
        RECT  4.795 1.515 5.185 1.715 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.105 -0.250 9.660 0.250 ;
        RECT  8.845 -0.250 9.105 0.405 ;
        RECT  8.025 -0.250 8.845 0.250 ;
        RECT  7.765 -0.250 8.025 0.405 ;
        RECT  6.455 -0.250 7.765 0.250 ;
        RECT  6.295 -0.250 6.455 0.625 ;
        RECT  5.095 -0.250 6.295 0.250 ;
        RECT  4.935 -0.250 5.095 0.690 ;
        RECT  4.065 -0.250 4.935 0.250 ;
        RECT  3.805 -0.250 4.065 0.875 ;
        RECT  1.790 -0.250 3.805 0.250 ;
        RECT  1.530 -0.250 1.790 0.405 ;
        RECT  0.385 -0.250 1.530 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.120 3.440 9.660 3.940 ;
        RECT  8.860 3.285 9.120 3.940 ;
        RECT  8.070 3.440 8.860 3.940 ;
        RECT  7.810 2.785 8.070 3.940 ;
        RECT  7.775 3.285 7.810 3.940 ;
        RECT  5.640 3.440 7.775 3.940 ;
        RECT  5.380 3.285 5.640 3.940 ;
        RECT  3.780 3.440 5.380 3.940 ;
        RECT  3.520 3.285 3.780 3.940 ;
        RECT  1.755 3.440 3.520 3.940 ;
        RECT  1.495 3.285 1.755 3.940 ;
        RECT  0.385 3.440 1.495 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.635 1.475 8.805 1.735 ;
        RECT  8.475 1.105 8.635 2.395 ;
        RECT  8.335 1.105 8.475 1.365 ;
        RECT  8.350 2.135 8.475 2.395 ;
        RECT  7.435 2.185 8.350 2.345 ;
        RECT  8.035 1.545 8.295 1.805 ;
        RECT  7.095 1.645 8.035 1.805 ;
        RECT  7.435 2.850 7.615 3.110 ;
        RECT  6.850 0.430 7.475 0.590 ;
        RECT  7.275 2.185 7.435 3.135 ;
        RECT  7.095 1.085 7.275 1.345 ;
        RECT  6.525 2.975 7.275 3.135 ;
        RECT  7.015 1.085 7.095 2.740 ;
        RECT  6.965 1.160 7.015 2.740 ;
        RECT  6.935 1.160 6.965 2.790 ;
        RECT  6.705 2.530 6.935 2.790 ;
        RECT  6.690 0.430 6.850 0.980 ;
        RECT  6.525 2.190 6.755 2.350 ;
        RECT  6.525 0.805 6.690 0.980 ;
        RECT  6.365 0.805 6.525 2.765 ;
        RECT  6.365 2.945 6.525 3.135 ;
        RECT  6.115 0.805 6.365 0.965 ;
        RECT  4.560 2.605 6.365 2.765 ;
        RECT  4.940 2.945 6.365 3.105 ;
        RECT  6.025 1.485 6.185 2.410 ;
        RECT  5.955 0.430 6.115 0.965 ;
        RECT  5.975 1.485 6.025 1.645 ;
        RECT  5.165 2.250 6.025 2.410 ;
        RECT  5.935 1.355 5.975 1.645 ;
        RECT  5.435 0.430 5.955 0.590 ;
        RECT  5.775 1.145 5.935 1.645 ;
        RECT  5.585 1.895 5.845 2.065 ;
        RECT  5.615 0.770 5.775 1.305 ;
        RECT  4.595 1.895 5.585 2.055 ;
        RECT  5.275 0.430 5.435 1.060 ;
        RECT  4.805 0.900 5.275 1.060 ;
        RECT  4.905 2.235 5.165 2.410 ;
        RECT  4.780 2.945 4.940 3.260 ;
        RECT  4.645 0.900 4.805 1.335 ;
        RECT  4.120 3.100 4.780 3.260 ;
        RECT  4.465 0.550 4.635 0.710 ;
        RECT  4.465 1.895 4.595 2.215 ;
        RECT  4.460 2.605 4.560 2.920 ;
        RECT  4.305 0.550 4.465 2.215 ;
        RECT  4.300 2.500 4.460 2.920 ;
        RECT  3.865 1.185 4.305 1.345 ;
        RECT  2.795 2.500 4.300 2.660 ;
        RECT  3.965 1.565 4.125 1.825 ;
        RECT  3.960 2.940 4.120 3.260 ;
        RECT  3.135 1.565 3.965 1.725 ;
        RECT  1.065 2.940 3.960 3.100 ;
        RECT  3.605 1.085 3.865 1.345 ;
        RECT  3.135 0.745 3.185 1.005 ;
        RECT  2.975 0.745 3.135 2.265 ;
        RECT  2.925 0.745 2.975 1.005 ;
        RECT  2.635 1.185 2.795 2.660 ;
        RECT  2.465 1.185 2.635 1.345 ;
        RECT  2.515 0.745 2.615 1.005 ;
        RECT  2.355 0.585 2.515 1.005 ;
        RECT  2.295 2.300 2.455 2.660 ;
        RECT  0.895 0.585 2.355 0.745 ;
        RECT  0.815 2.500 2.295 2.660 ;
        RECT  1.595 1.910 1.855 2.170 ;
        RECT  1.510 1.910 1.595 2.070 ;
        RECT  1.350 1.165 1.510 2.070 ;
        RECT  0.765 1.165 1.350 1.325 ;
        RECT  0.805 2.940 1.065 3.200 ;
        RECT  0.685 0.430 0.895 0.745 ;
        RECT  0.765 1.960 0.815 2.220 ;
        RECT  0.555 2.500 0.815 2.760 ;
        RECT  0.605 1.035 0.765 2.220 ;
        RECT  0.635 0.430 0.685 0.690 ;
        RECT  0.555 1.960 0.605 2.220 ;
    END
END EDFFXL

MACRO DFFTRX4
    CLASS CORE ;
    FOREIGN DFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.435 0.405 1.995 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 1.290 9.535 1.990 ;
        RECT  9.320 1.290 9.380 3.215 ;
        RECT  9.120 1.035 9.320 3.215 ;
        RECT  9.015 1.035 9.120 1.295 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.400 0.945 10.455 2.995 ;
        RECT  10.165 0.695 10.400 3.215 ;
        RECT  10.140 0.695 10.165 1.295 ;
        RECT  10.140 2.275 10.165 3.215 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.685 1.290 1.035 1.940 ;
        RECT  0.585 1.290 0.685 1.765 ;
        END
        ANTENNAGATEAREA     0.2392 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.380 1.610 ;
        END
        ANTENNAGATEAREA     0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.910 -0.250 11.040 0.250 ;
        RECT  10.650 -0.250 10.910 1.130 ;
        RECT  9.820 -0.250 10.650 0.250 ;
        RECT  9.560 -0.250 9.820 0.405 ;
        RECT  8.710 -0.250 9.560 0.250 ;
        RECT  8.450 -0.250 8.710 0.405 ;
        RECT  7.635 -0.250 8.450 0.250 ;
        RECT  7.375 -0.250 7.635 1.295 ;
        RECT  5.005 -0.250 7.375 0.250 ;
        RECT  4.745 -0.250 5.005 0.575 ;
        RECT  4.385 -0.250 4.745 0.250 ;
        RECT  4.125 -0.250 4.385 0.655 ;
        RECT  2.425 -0.250 4.125 0.250 ;
        RECT  2.165 -0.250 2.425 0.405 ;
        RECT  0.385 -0.250 2.165 0.250 ;
        RECT  0.125 -0.250 0.385 1.115 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.910 3.440 11.040 3.940 ;
        RECT  10.650 2.220 10.910 3.940 ;
        RECT  9.890 3.440 10.650 3.940 ;
        RECT  9.630 2.275 9.890 3.940 ;
        RECT  8.870 3.440 9.630 3.940 ;
        RECT  8.610 2.260 8.870 3.940 ;
        RECT  7.780 3.440 8.610 3.940 ;
        RECT  7.520 3.285 7.780 3.940 ;
        RECT  5.260 3.440 7.520 3.940 ;
        RECT  5.000 2.640 5.260 3.940 ;
        RECT  4.240 3.440 5.000 3.940 ;
        RECT  3.980 2.725 4.240 3.940 ;
        RECT  2.770 3.440 3.980 3.940 ;
        RECT  2.510 3.285 2.770 3.940 ;
        RECT  0.785 3.440 2.510 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.955 1.535 9.985 1.795 ;
        RECT  9.795 0.690 9.955 1.795 ;
        RECT  8.835 0.690 9.795 0.850 ;
        RECT  8.675 0.690 8.835 1.145 ;
        RECT  8.255 0.985 8.675 1.145 ;
        RECT  8.255 1.955 8.355 2.555 ;
        RECT  8.095 0.985 8.255 2.555 ;
        RECT  7.925 2.735 8.185 2.995 ;
        RECT  7.915 0.985 8.095 1.245 ;
        RECT  7.225 1.585 8.095 1.915 ;
        RECT  6.630 2.735 7.925 2.895 ;
        RECT  6.885 0.470 7.045 2.405 ;
        RECT  5.345 0.470 6.885 0.630 ;
        RECT  6.845 2.140 6.885 2.405 ;
        RECT  6.630 0.985 6.705 1.245 ;
        RECT  6.470 0.815 6.630 3.020 ;
        RECT  5.685 0.815 6.470 0.975 ;
        RECT  5.660 2.860 6.470 3.020 ;
        RECT  6.170 1.160 6.245 1.320 ;
        RECT  5.985 1.160 6.170 2.645 ;
        RECT  5.085 1.485 5.985 1.650 ;
        RECT  5.910 2.045 5.985 2.645 ;
        RECT  5.525 0.815 5.685 1.300 ;
        RECT  5.500 2.045 5.660 3.020 ;
        RECT  5.400 2.045 5.500 2.305 ;
        RECT  5.185 0.470 5.345 0.995 ;
        RECT  3.835 0.835 5.185 0.995 ;
        RECT  4.925 1.485 5.085 2.425 ;
        RECT  4.785 1.485 4.925 1.645 ;
        RECT  4.750 2.265 4.925 2.425 ;
        RECT  4.525 1.175 4.785 1.645 ;
        RECT  4.490 2.265 4.750 2.865 ;
        RECT  4.460 1.825 4.720 2.085 ;
        RECT  3.950 1.485 4.525 1.645 ;
        RECT  4.290 1.925 4.460 2.085 ;
        RECT  4.130 1.925 4.290 2.330 ;
        RECT  3.610 2.165 4.130 2.330 ;
        RECT  3.790 1.485 3.950 1.985 ;
        RECT  3.690 0.695 3.835 0.995 ;
        RECT  3.675 0.590 3.690 0.995 ;
        RECT  3.430 0.590 3.675 0.855 ;
        RECT  3.450 1.650 3.610 2.845 ;
        RECT  3.435 1.650 3.450 1.810 ;
        RECT  3.350 2.685 3.450 2.845 ;
        RECT  3.275 1.035 3.435 1.810 ;
        RECT  3.095 0.640 3.430 0.855 ;
        RECT  3.090 2.685 3.350 2.945 ;
        RECT  3.095 2.005 3.270 2.265 ;
        RECT  2.935 0.575 3.095 2.505 ;
        RECT  1.850 2.785 3.090 2.945 ;
        RECT  2.755 0.575 2.935 0.735 ;
        RECT  2.060 2.345 2.935 2.505 ;
        RECT  2.595 0.950 2.755 2.165 ;
        RECT  2.025 0.950 2.595 1.110 ;
        RECT  2.050 2.005 2.595 2.165 ;
        RECT  1.900 2.345 2.060 2.605 ;
        RECT  1.925 0.850 2.025 1.110 ;
        RECT  1.765 0.430 1.925 1.110 ;
        RECT  1.720 2.785 1.850 3.075 ;
        RECT  1.515 0.430 1.765 0.590 ;
        RECT  1.560 1.490 1.720 3.075 ;
        RECT  1.515 1.490 1.560 1.650 ;
        RECT  1.355 1.035 1.515 1.650 ;
        RECT  1.255 1.035 1.355 1.295 ;
        RECT  1.080 2.135 1.340 3.075 ;
        RECT  0.385 2.315 1.080 2.475 ;
        RECT  0.125 2.315 0.385 2.575 ;
    END
END DFFTRX4

MACRO DFFTRX2
    CLASS CORE ;
    FOREIGN DFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 1.285 1.380 1.545 ;
        RECT  1.045 1.285 1.320 1.990 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.075 1.290 7.235 1.580 ;
        RECT  7.035 2.160 7.135 3.100 ;
        RECT  7.035 1.000 7.075 1.580 ;
        RECT  6.875 1.000 7.035 3.100 ;
        RECT  6.815 1.000 6.875 1.260 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.995 0.695 8.155 3.125 ;
        RECT  7.895 0.695 7.995 1.295 ;
        RECT  7.895 2.185 7.995 3.125 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.845 1.855 ;
        END
        ANTENNAGATEAREA     0.1222 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.760 1.290 2.175 1.610 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.615 -0.250 8.280 0.250 ;
        RECT  7.355 -0.250 7.615 0.405 ;
        RECT  5.995 -0.250 7.355 0.250 ;
        RECT  5.735 -0.250 5.995 1.225 ;
        RECT  3.870 -0.250 5.735 0.250 ;
        RECT  3.610 -0.250 3.870 0.630 ;
        RECT  2.460 -0.250 3.610 0.250 ;
        RECT  2.200 -0.250 2.460 0.405 ;
        RECT  1.440 -0.250 2.200 0.250 ;
        RECT  1.180 -0.250 1.440 0.405 ;
        RECT  0.000 -0.250 1.180 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.645 3.440 8.280 3.940 ;
        RECT  7.385 2.155 7.645 3.940 ;
        RECT  5.995 3.440 7.385 3.940 ;
        RECT  5.945 3.285 5.995 3.940 ;
        RECT  5.785 2.895 5.945 3.940 ;
        RECT  5.735 3.285 5.785 3.940 ;
        RECT  3.860 3.440 5.735 3.940 ;
        RECT  3.600 2.405 3.860 3.940 ;
        RECT  2.310 3.440 3.600 3.940 ;
        RECT  2.050 3.285 2.310 3.940 ;
        RECT  1.450 3.440 2.050 3.940 ;
        RECT  1.190 3.285 1.450 3.940 ;
        RECT  0.000 3.440 1.190 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.715 1.535 7.815 1.795 ;
        RECT  7.555 0.615 7.715 1.795 ;
        RECT  6.565 0.615 7.555 0.775 ;
        RECT  6.500 2.025 6.600 2.285 ;
        RECT  6.500 0.615 6.565 1.245 ;
        RECT  6.405 0.615 6.500 2.285 ;
        RECT  6.150 2.475 6.410 2.735 ;
        RECT  6.340 0.985 6.405 2.285 ;
        RECT  6.305 0.985 6.340 1.915 ;
        RECT  5.585 1.655 6.305 1.915 ;
        RECT  5.575 2.555 6.150 2.715 ;
        RECT  5.415 2.555 5.575 2.820 ;
        RECT  4.945 2.660 5.415 2.820 ;
        RECT  5.245 0.605 5.405 1.595 ;
        RECT  4.215 0.605 5.245 0.765 ;
        RECT  5.235 1.435 5.245 1.595 ;
        RECT  5.075 1.435 5.235 2.480 ;
        RECT  4.905 0.985 5.065 1.245 ;
        RECT  4.895 2.660 4.945 3.005 ;
        RECT  4.895 1.085 4.905 1.245 ;
        RECT  4.735 1.085 4.895 3.005 ;
        RECT  4.685 2.745 4.735 3.005 ;
        RECT  4.435 0.945 4.555 2.500 ;
        RECT  4.395 0.945 4.435 2.940 ;
        RECT  3.955 1.360 4.395 1.620 ;
        RECT  4.175 2.340 4.395 2.940 ;
        RECT  4.055 0.605 4.215 0.970 ;
        RECT  3.335 1.835 4.215 2.095 ;
        RECT  2.855 0.810 4.055 0.970 ;
        RECT  3.695 1.355 3.955 1.620 ;
        RECT  3.175 1.210 3.335 2.885 ;
        RECT  3.055 1.210 3.175 1.470 ;
        RECT  2.895 2.725 3.175 2.885 ;
        RECT  2.855 1.650 2.995 1.910 ;
        RECT  2.635 2.725 2.895 3.105 ;
        RECT  2.855 2.265 2.890 2.425 ;
        RECT  2.695 0.705 2.855 2.425 ;
        RECT  0.680 2.265 2.695 2.425 ;
        RECT  0.390 2.945 2.635 3.105 ;
        RECT  2.355 0.585 2.515 2.085 ;
        RECT  1.950 0.585 2.355 0.745 ;
        RECT  1.620 1.925 2.355 2.085 ;
        RECT  1.690 0.465 1.950 0.745 ;
        RECT  0.640 2.605 1.880 2.765 ;
        RECT  0.755 0.585 1.690 0.745 ;
        RECT  0.595 0.465 0.755 0.745 ;
        RECT  0.520 2.075 0.680 2.425 ;
        RECT  0.330 0.465 0.595 0.625 ;
        RECT  0.290 0.905 0.390 1.165 ;
        RECT  0.290 2.635 0.390 3.105 ;
        RECT  0.130 0.905 0.290 3.105 ;
    END
END DFFTRX2

MACRO DFFTRX1
    CLASS CORE ;
    FOREIGN DFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.440 1.265 1.715 1.715 ;
        END
        ANTENNAGATEAREA     0.0481 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.690 1.140 6.835 2.715 ;
        RECT  6.675 1.035 6.690 2.715 ;
        RECT  6.565 1.035 6.675 1.580 ;
        RECT  6.660 2.555 6.675 2.715 ;
        RECT  6.400 2.555 6.660 3.215 ;
        RECT  6.530 1.035 6.565 1.300 ;
        END
        ANTENNADIFFAREA     0.3472 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.690 1.105 7.695 2.995 ;
        RECT  7.530 0.995 7.690 3.215 ;
        RECT  7.485 0.995 7.530 1.365 ;
        RECT  7.485 2.335 7.530 3.215 ;
        RECT  7.430 0.995 7.485 1.255 ;
        RECT  7.480 2.585 7.485 3.215 ;
        RECT  7.430 2.615 7.480 3.215 ;
        END
        ANTENNADIFFAREA     0.3468 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.700 1.255 1.990 ;
        RECT  0.810 1.705 1.045 1.965 ;
        END
        ANTENNAGATEAREA     0.0676 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.165 1.265 2.175 1.580 ;
        RECT  1.900 1.265 2.165 1.715 ;
        END
        ANTENNAGATEAREA     0.0468 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.215 -0.250 7.820 0.250 ;
        RECT  6.955 -0.250 7.215 0.405 ;
        RECT  5.790 -0.250 6.955 0.250 ;
        RECT  5.530 -0.250 5.790 0.405 ;
        RECT  4.150 -0.250 5.530 0.250 ;
        RECT  3.890 -0.250 4.150 1.150 ;
        RECT  2.460 -0.250 3.890 0.250 ;
        RECT  2.200 -0.250 2.460 0.405 ;
        RECT  1.440 -0.250 2.200 0.250 ;
        RECT  1.180 -0.250 1.440 0.405 ;
        RECT  0.000 -0.250 1.180 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.170 3.440 7.820 3.940 ;
        RECT  6.910 2.925 7.170 3.940 ;
        RECT  5.990 3.440 6.910 3.940 ;
        RECT  5.730 2.865 5.990 3.940 ;
        RECT  3.805 3.440 5.730 3.940 ;
        RECT  3.545 2.650 3.805 3.940 ;
        RECT  2.310 3.440 3.545 3.940 ;
        RECT  2.050 3.285 2.310 3.940 ;
        RECT  1.450 3.440 2.050 3.940 ;
        RECT  1.190 3.285 1.450 3.940 ;
        RECT  0.000 3.440 1.190 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.175 1.725 7.350 1.985 ;
        RECT  7.015 0.685 7.175 1.985 ;
        RECT  6.335 0.685 7.015 0.845 ;
        RECT  6.335 2.105 6.495 2.365 ;
        RECT  6.175 0.495 6.335 2.365 ;
        RECT  6.040 0.495 6.175 0.755 ;
        RECT  5.560 1.125 6.175 1.285 ;
        RECT  5.830 1.465 5.990 2.615 ;
        RECT  5.100 2.455 5.830 2.615 ;
        RECT  5.560 1.945 5.610 2.205 ;
        RECT  5.400 1.125 5.560 2.205 ;
        RECT  5.350 1.945 5.400 2.205 ;
        RECT  5.040 2.960 5.300 3.220 ;
        RECT  5.100 0.490 5.190 0.650 ;
        RECT  4.940 0.490 5.100 2.760 ;
        RECT  4.175 3.010 5.040 3.170 ;
        RECT  4.930 0.490 4.940 0.650 ;
        RECT  4.840 2.500 4.940 2.760 ;
        RECT  4.515 1.530 4.750 1.790 ;
        RECT  4.355 1.405 4.515 2.770 ;
        RECT  3.850 1.405 4.355 1.665 ;
        RECT  4.015 1.865 4.175 3.170 ;
        RECT  3.670 1.865 4.015 2.025 ;
        RECT  3.330 2.210 3.835 2.470 ;
        RECT  3.510 0.790 3.670 2.025 ;
        RECT  2.970 0.790 3.510 0.950 ;
        RECT  3.170 1.210 3.330 2.740 ;
        RECT  3.050 1.210 3.170 1.475 ;
        RECT  2.895 2.580 3.170 2.740 ;
        RECT  2.870 1.660 2.990 1.920 ;
        RECT  2.870 0.630 2.970 0.950 ;
        RECT  2.845 2.580 2.895 2.955 ;
        RECT  2.870 2.235 2.890 2.395 ;
        RECT  2.710 0.630 2.870 2.395 ;
        RECT  2.735 2.580 2.845 3.105 ;
        RECT  2.635 2.695 2.735 3.105 ;
        RECT  0.470 2.235 2.710 2.395 ;
        RECT  0.340 2.945 2.635 3.105 ;
        RECT  2.370 0.885 2.530 2.055 ;
        RECT  1.950 0.885 2.370 1.045 ;
        RECT  2.350 1.745 2.370 2.055 ;
        RECT  1.620 1.895 2.350 2.055 ;
        RECT  1.790 0.435 1.950 1.045 ;
        RECT  0.640 2.605 1.880 2.765 ;
        RECT  1.690 0.435 1.790 0.745 ;
        RECT  0.590 0.585 1.690 0.745 ;
        RECT  0.330 0.565 0.590 0.825 ;
        RECT  0.290 1.005 0.390 1.265 ;
        RECT  0.290 2.555 0.340 3.105 ;
        RECT  0.130 1.005 0.290 3.105 ;
    END
END DFFTRX1

MACRO DFFTRXL
    CLASS CORE ;
    FOREIGN DFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 1.265 1.720 1.665 ;
        RECT  1.300 1.265 1.435 1.505 ;
        END
        ANTENNAGATEAREA     0.0403 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.765 1.135 6.925 2.945 ;
        RECT  6.660 1.135 6.765 1.295 ;
        RECT  6.545 2.785 6.765 2.945 ;
        RECT  6.400 1.035 6.660 1.295 ;
        RECT  6.315 2.785 6.545 3.195 ;
        RECT  6.105 2.930 6.315 3.220 ;
        END
        ANTENNADIFFAREA     0.2142 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.635 1.355 7.695 2.995 ;
        RECT  7.630 1.355 7.635 3.195 ;
        RECT  7.470 1.035 7.630 3.195 ;
        RECT  7.465 2.685 7.470 3.195 ;
        RECT  7.375 2.935 7.465 3.195 ;
        END
        ANTENNADIFFAREA     0.2164 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.070 1.700 1.255 1.990 ;
        RECT  1.045 1.685 1.070 1.990 ;
        RECT  0.810 1.685 1.045 1.945 ;
        END
        ANTENNAGATEAREA     0.0468 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.265 2.280 1.565 ;
        RECT  1.900 1.265 2.175 1.635 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.240 -0.250 7.820 0.250 ;
        RECT  6.980 -0.250 7.240 0.405 ;
        RECT  6.045 -0.250 6.980 0.250 ;
        RECT  5.785 -0.250 6.045 0.405 ;
        RECT  4.250 -0.250 5.785 0.250 ;
        RECT  3.990 -0.250 4.250 1.150 ;
        RECT  2.380 -0.250 3.990 0.250 ;
        RECT  2.120 -0.250 2.380 0.405 ;
        RECT  1.590 -0.250 2.120 0.250 ;
        RECT  1.330 -0.250 1.590 0.405 ;
        RECT  0.000 -0.250 1.330 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.090 3.440 7.820 3.940 ;
        RECT  6.830 3.125 7.090 3.940 ;
        RECT  5.840 3.440 6.830 3.940 ;
        RECT  5.580 2.870 5.840 3.940 ;
        RECT  3.775 3.440 5.580 3.940 ;
        RECT  3.515 2.505 3.775 3.940 ;
        RECT  2.310 3.440 3.515 3.940 ;
        RECT  2.050 3.285 2.310 3.940 ;
        RECT  1.450 3.440 2.050 3.940 ;
        RECT  1.190 3.285 1.450 3.940 ;
        RECT  0.000 3.440 1.190 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.130 0.620 7.290 1.760 ;
        RECT  6.660 0.620 7.130 0.780 ;
        RECT  6.400 0.520 6.660 0.780 ;
        RECT  6.420 1.480 6.580 2.605 ;
        RECT  6.000 1.480 6.420 1.640 ;
        RECT  6.165 2.445 6.420 2.605 ;
        RECT  6.000 0.615 6.400 0.780 ;
        RECT  6.080 1.985 6.240 2.245 ;
        RECT  5.295 1.985 6.080 2.145 ;
        RECT  5.840 0.615 6.000 1.640 ;
        RECT  5.720 1.310 5.840 1.570 ;
        RECT  5.295 0.455 5.400 0.715 ;
        RECT  5.040 2.865 5.300 3.125 ;
        RECT  5.140 0.455 5.295 2.145 ;
        RECT  5.135 0.505 5.140 2.145 ;
        RECT  5.100 1.985 5.135 2.145 ;
        RECT  4.940 1.985 5.100 2.685 ;
        RECT  4.175 2.865 5.040 3.025 ;
        RECT  4.840 2.425 4.940 2.685 ;
        RECT  4.720 0.940 4.820 1.200 ;
        RECT  4.560 0.940 4.720 1.520 ;
        RECT  4.515 1.360 4.560 1.520 ;
        RECT  4.355 1.360 4.515 2.685 ;
        RECT  3.880 1.360 4.355 1.520 ;
        RECT  4.015 1.700 4.175 3.025 ;
        RECT  3.700 1.700 4.015 1.860 ;
        RECT  3.360 2.040 3.835 2.300 ;
        RECT  3.540 0.680 3.700 1.860 ;
        RECT  3.005 0.680 3.540 0.840 ;
        RECT  3.335 1.020 3.360 2.300 ;
        RECT  3.200 1.020 3.335 2.840 ;
        RECT  3.160 1.020 3.200 1.280 ;
        RECT  3.175 2.090 3.200 2.840 ;
        RECT  2.895 2.680 3.175 2.840 ;
        RECT  2.965 1.415 3.020 1.675 ;
        RECT  2.965 0.515 3.005 0.840 ;
        RECT  2.805 0.515 2.965 2.445 ;
        RECT  2.795 2.680 2.895 2.955 ;
        RECT  2.745 0.515 2.805 0.775 ;
        RECT  2.630 2.185 2.805 2.445 ;
        RECT  2.635 2.680 2.795 3.105 ;
        RECT  0.290 2.945 2.635 3.105 ;
        RECT  0.710 2.235 2.630 2.395 ;
        RECT  2.460 0.925 2.620 2.005 ;
        RECT  0.750 0.925 2.460 1.085 ;
        RECT  2.380 1.745 2.460 2.005 ;
        RECT  1.880 1.845 2.380 2.005 ;
        RECT  1.620 1.845 1.880 2.055 ;
        RECT  0.565 2.605 1.880 2.765 ;
        RECT  0.590 0.695 0.750 1.085 ;
        RECT  0.550 2.165 0.710 2.425 ;
        RECT  0.330 0.595 0.590 0.855 ;
        RECT  0.290 1.035 0.390 1.295 ;
        RECT  0.290 1.955 0.340 2.215 ;
        RECT  0.130 1.035 0.290 3.105 ;
    END
END DFFTRXL

MACRO DFFNSRX4
    CLASS CORE ;
    FOREIGN DFFNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.665 2.930 11.835 3.220 ;
        RECT  11.500 2.520 11.665 3.220 ;
        RECT  11.380 2.520 11.500 2.810 ;
        END
        ANTENNAGATEAREA     0.3250 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.700 4.015 1.990 ;
        RECT  3.805 1.680 4.005 1.990 ;
        RECT  3.460 1.680 3.805 1.985 ;
        END
        ANTENNAGATEAREA     0.1027 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.995 0.595 14.155 2.320 ;
        RECT  12.495 0.595 13.995 0.755 ;
        RECT  13.210 2.160 13.995 2.320 ;
        RECT  13.210 2.520 13.215 3.220 ;
        RECT  13.005 2.160 13.210 3.220 ;
        RECT  12.940 2.160 13.005 3.100 ;
        RECT  12.235 0.595 12.495 1.195 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.860 1.290 15.055 1.990 ;
        RECT  14.845 1.085 14.860 1.990 ;
        RECT  14.495 1.085 14.845 2.745 ;
        RECT  14.385 0.645 14.495 2.745 ;
        RECT  14.335 0.645 14.385 1.245 ;
        RECT  14.220 2.505 14.385 2.745 ;
        RECT  13.960 2.505 14.220 3.105 ;
        RECT  13.925 2.745 13.960 3.000 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 1.405 0.585 1.665 ;
        RECT  0.125 1.285 0.445 1.665 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.710 1.695 3.180 1.990 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.055 -0.250 15.180 0.250 ;
        RECT  14.795 -0.250 15.055 0.795 ;
        RECT  13.995 -0.250 14.795 0.250 ;
        RECT  13.735 -0.250 13.995 0.405 ;
        RECT  13.045 -0.250 13.735 0.250 ;
        RECT  12.785 -0.250 13.045 0.405 ;
        RECT  11.985 -0.250 12.785 0.250 ;
        RECT  11.725 -0.250 11.985 1.165 ;
        RECT  10.925 -0.250 11.725 0.250 ;
        RECT  10.665 -0.250 10.925 1.135 ;
        RECT  3.485 -0.250 10.665 0.250 ;
        RECT  3.225 -0.250 3.485 0.405 ;
        RECT  2.315 -0.250 3.225 0.250 ;
        RECT  2.055 -0.250 2.315 0.405 ;
        RECT  0.475 -0.250 2.055 0.250 ;
        RECT  0.215 -0.250 0.475 1.075 ;
        RECT  0.000 -0.250 0.215 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.745 3.440 15.180 3.940 ;
        RECT  14.485 2.955 14.745 3.940 ;
        RECT  13.710 3.440 14.485 3.940 ;
        RECT  13.450 2.600 13.710 3.940 ;
        RECT  12.665 3.440 13.450 3.940 ;
        RECT  12.405 2.445 12.665 3.940 ;
        RECT  9.440 3.440 12.405 3.940 ;
        RECT  8.840 3.285 9.440 3.940 ;
        RECT  6.140 3.440 8.840 3.940 ;
        RECT  5.880 3.105 6.140 3.940 ;
        RECT  4.430 3.440 5.880 3.940 ;
        RECT  3.830 3.055 4.430 3.940 ;
        RECT  2.245 3.440 3.830 3.940 ;
        RECT  1.985 3.285 2.245 3.940 ;
        RECT  0.430 3.440 1.985 3.940 ;
        RECT  0.170 2.195 0.430 3.940 ;
        RECT  0.000 3.440 0.170 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.640 0.955 13.800 1.980 ;
        RECT  13.185 0.955 13.640 1.115 ;
        RECT  12.610 1.820 13.640 1.980 ;
        RECT  12.225 1.470 13.345 1.630 ;
        RECT  12.450 1.820 12.610 2.265 ;
        RECT  12.155 2.105 12.450 2.265 ;
        RECT  12.065 1.470 12.225 1.905 ;
        RECT  11.895 2.105 12.155 2.740 ;
        RECT  10.100 1.745 12.065 1.905 ;
        RECT  11.000 2.105 11.895 2.265 ;
        RECT  11.215 0.495 11.475 1.565 ;
        RECT  10.480 1.405 11.215 1.565 ;
        RECT  10.940 2.890 11.200 3.150 ;
        RECT  10.740 2.085 11.000 2.345 ;
        RECT  6.690 2.945 10.940 3.105 ;
        RECT  10.320 0.470 10.480 1.565 ;
        RECT  10.310 2.500 10.470 2.765 ;
        RECT  6.520 0.470 10.320 0.630 ;
        RECT  7.095 2.605 10.310 2.765 ;
        RECT  10.100 2.245 10.150 2.405 ;
        RECT  9.940 0.815 10.100 2.405 ;
        RECT  8.375 0.815 9.940 0.975 ;
        RECT  7.810 2.245 9.940 2.405 ;
        RECT  9.420 1.160 9.680 1.455 ;
        RECT  8.060 1.160 9.420 1.320 ;
        RECT  7.630 1.505 9.225 1.665 ;
        RECT  7.900 0.820 8.060 1.320 ;
        RECT  7.005 0.820 7.900 0.980 ;
        RECT  7.470 1.160 7.630 2.245 ;
        RECT  7.195 1.160 7.470 1.320 ;
        RECT  6.335 2.085 7.470 2.245 ;
        RECT  7.005 1.560 7.290 1.830 ;
        RECT  6.935 2.425 7.095 2.765 ;
        RECT  6.845 0.820 7.005 1.830 ;
        RECT  4.945 2.425 6.935 2.585 ;
        RECT  6.180 0.940 6.845 1.100 ;
        RECT  6.530 2.765 6.690 3.105 ;
        RECT  6.430 2.765 6.530 2.940 ;
        RECT  6.360 0.470 6.520 0.755 ;
        RECT  5.590 2.765 6.430 2.925 ;
        RECT  6.175 1.335 6.335 2.245 ;
        RECT  6.020 0.585 6.180 1.100 ;
        RECT  5.840 1.335 6.175 1.495 ;
        RECT  4.780 2.085 6.175 2.245 ;
        RECT  2.895 0.585 6.020 0.745 ;
        RECT  5.680 0.965 5.840 1.495 ;
        RECT  5.580 0.965 5.680 1.225 ;
        RECT  5.320 2.765 5.590 2.940 ;
        RECT  4.895 1.065 5.580 1.225 ;
        RECT  4.785 2.425 4.945 2.870 ;
        RECT  4.630 0.925 4.895 1.225 ;
        RECT  3.420 2.710 4.785 2.870 ;
        RECT  2.115 0.925 4.630 1.085 ;
        RECT  4.360 1.680 4.600 1.940 ;
        RECT  4.360 2.365 4.520 2.525 ;
        RECT  4.200 1.275 4.360 2.525 ;
        RECT  3.790 1.275 4.200 1.435 ;
        RECT  3.260 2.170 3.420 2.910 ;
        RECT  2.495 2.170 3.260 2.330 ;
        RECT  3.080 3.100 3.185 3.260 ;
        RECT  2.920 2.510 3.080 3.260 ;
        RECT  1.450 2.510 2.920 2.670 ;
        RECT  2.635 0.525 2.895 0.745 ;
        RECT  2.495 1.275 2.885 1.435 ;
        RECT  2.580 2.850 2.740 3.110 ;
        RECT  0.930 0.585 2.635 0.745 ;
        RECT  0.775 2.885 2.580 3.045 ;
        RECT  2.335 1.275 2.495 2.330 ;
        RECT  1.795 1.695 2.335 1.855 ;
        RECT  1.955 0.925 2.115 1.425 ;
        RECT  1.635 1.650 1.795 1.910 ;
        RECT  1.425 2.290 1.450 2.670 ;
        RECT  1.265 0.935 1.425 2.670 ;
        RECT  1.115 0.935 1.265 1.095 ;
        RECT  1.110 2.070 1.265 2.670 ;
        RECT  0.930 1.355 1.085 1.615 ;
        RECT  0.775 0.585 0.930 2.005 ;
        RECT  0.770 0.585 0.775 3.045 ;
        RECT  0.615 1.845 0.770 3.045 ;
    END
END DFFNSRX4

MACRO DFFNSRX2
    CLASS CORE ;
    FOREIGN DFFNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.405 2.930 8.615 3.220 ;
        RECT  8.110 2.960 8.405 3.220 ;
        END
        ANTENNAGATEAREA     0.1703 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.680 3.720 1.985 ;
        RECT  3.345 1.680 3.555 1.990 ;
        RECT  3.275 1.680 3.345 1.985 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.245 0.585 10.455 2.420 ;
        RECT  9.435 0.585 10.245 0.745 ;
        RECT  9.975 2.260 10.245 2.420 ;
        RECT  9.715 2.260 9.975 2.520 ;
        RECT  9.175 0.585 9.435 1.235 ;
        END
        ANTENNADIFFAREA     0.6007 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.655 0.645 10.915 3.025 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.520 0.370 1.990 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.625 1.695 3.095 1.990 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.375 -0.250 11.040 0.250 ;
        RECT  10.115 -0.250 10.375 0.405 ;
        RECT  8.925 -0.250 10.115 0.250 ;
        RECT  8.665 -0.250 8.925 1.165 ;
        RECT  3.345 -0.250 8.665 0.250 ;
        RECT  3.085 -0.250 3.345 0.405 ;
        RECT  2.185 -0.250 3.085 0.250 ;
        RECT  1.925 -0.250 2.185 0.405 ;
        RECT  0.385 -0.250 1.925 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 3.440 11.040 3.940 ;
        RECT  10.145 2.935 10.405 3.940 ;
        RECT  9.465 3.440 10.145 3.940 ;
        RECT  9.205 2.275 9.465 3.940 ;
        RECT  6.725 3.440 9.205 3.940 ;
        RECT  6.465 3.115 6.725 3.940 ;
        RECT  5.305 3.440 6.465 3.940 ;
        RECT  5.145 2.825 5.305 3.940 ;
        RECT  4.185 3.440 5.145 3.940 ;
        RECT  3.585 3.055 4.185 3.940 ;
        RECT  2.005 3.440 3.585 3.940 ;
        RECT  1.745 3.285 2.005 3.940 ;
        RECT  0.385 3.440 1.745 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.905 0.965 10.065 2.005 ;
        RECT  9.685 0.965 9.905 1.125 ;
        RECT  8.815 1.845 9.905 2.005 ;
        RECT  8.980 1.455 9.495 1.615 ;
        RECT  8.820 1.350 8.980 1.615 ;
        RECT  7.800 1.350 8.820 1.510 ;
        RECT  8.555 1.845 8.815 2.565 ;
        RECT  8.045 1.845 8.555 2.005 ;
        RECT  8.075 0.470 8.335 1.075 ;
        RECT  7.825 2.405 8.085 2.665 ;
        RECT  7.995 0.470 8.075 0.630 ;
        RECT  7.785 1.745 8.045 2.005 ;
        RECT  7.835 0.430 7.995 0.630 ;
        RECT  7.215 0.430 7.835 0.590 ;
        RECT  7.800 2.505 7.825 2.665 ;
        RECT  7.640 1.155 7.800 1.510 ;
        RECT  7.640 2.505 7.800 2.935 ;
        RECT  7.395 0.775 7.655 0.970 ;
        RECT  7.120 1.155 7.640 1.315 ;
        RECT  5.675 2.775 7.640 2.935 ;
        RECT  7.300 1.635 7.460 2.595 ;
        RECT  6.780 0.810 7.395 0.970 ;
        RECT  6.015 2.435 7.300 2.595 ;
        RECT  7.055 0.430 7.215 0.630 ;
        RECT  6.960 1.155 7.120 2.235 ;
        RECT  5.280 0.470 7.055 0.630 ;
        RECT  6.745 2.075 6.960 2.235 ;
        RECT  6.620 0.810 6.780 1.885 ;
        RECT  5.625 0.810 6.620 0.970 ;
        RECT  6.535 1.625 6.620 1.885 ;
        RECT  6.355 2.075 6.495 2.235 ;
        RECT  6.355 1.150 6.410 1.310 ;
        RECT  6.195 1.150 6.355 2.235 ;
        RECT  5.810 1.150 6.195 1.445 ;
        RECT  5.855 1.975 6.015 2.595 ;
        RECT  4.425 1.975 5.855 2.135 ;
        RECT  4.600 1.285 5.810 1.445 ;
        RECT  5.515 2.315 5.675 2.935 ;
        RECT  5.465 0.810 5.625 1.100 ;
        RECT  4.765 2.315 5.515 2.475 ;
        RECT  4.940 0.940 5.465 1.100 ;
        RECT  5.120 0.470 5.280 0.755 ;
        RECT  4.780 0.545 4.940 1.100 ;
        RECT  3.690 0.545 4.780 0.705 ;
        RECT  4.605 2.315 4.765 2.920 ;
        RECT  4.085 1.635 4.645 1.795 ;
        RECT  4.440 0.890 4.600 1.445 ;
        RECT  4.390 0.890 4.440 1.145 ;
        RECT  4.265 1.975 4.425 2.755 ;
        RECT  2.025 0.925 4.390 1.085 ;
        RECT  3.215 2.595 4.265 2.755 ;
        RECT  3.925 1.265 4.085 2.375 ;
        RECT  3.670 1.265 3.925 1.425 ;
        RECT  3.575 2.215 3.925 2.375 ;
        RECT  3.530 0.545 3.690 0.745 ;
        RECT  2.785 0.585 3.530 0.745 ;
        RECT  3.055 2.170 3.215 2.910 ;
        RECT  2.395 2.170 3.055 2.330 ;
        RECT  2.875 3.100 2.975 3.260 ;
        RECT  2.715 2.510 2.875 3.260 ;
        RECT  2.525 0.445 2.785 0.745 ;
        RECT  2.365 1.275 2.775 1.435 ;
        RECT  1.265 2.510 2.715 2.670 ;
        RECT  2.375 2.850 2.535 3.110 ;
        RECT  0.820 0.585 2.525 0.745 ;
        RECT  2.365 2.015 2.395 2.330 ;
        RECT  1.465 2.850 2.375 3.010 ;
        RECT  2.205 1.275 2.365 2.330 ;
        RECT  2.135 1.645 2.205 2.330 ;
        RECT  1.555 1.645 2.135 1.805 ;
        RECT  1.865 0.925 2.025 1.425 ;
        RECT  1.395 1.645 1.555 1.910 ;
        RECT  1.205 2.850 1.465 3.120 ;
        RECT  1.215 0.945 1.395 1.205 ;
        RECT  1.215 2.270 1.265 2.670 ;
        RECT  1.055 0.945 1.215 2.670 ;
        RECT  0.820 2.850 1.205 3.010 ;
        RECT  1.005 2.270 1.055 2.530 ;
        RECT  0.820 1.320 0.875 1.580 ;
        RECT  0.660 0.585 0.820 3.010 ;
    END
END DFFNSRX2

MACRO DFFNSRX1
    CLASS CORE ;
    FOREIGN DFFNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.750 2.865 8.155 3.220 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.700 3.885 1.960 ;
        RECT  3.525 1.290 3.555 1.960 ;
        RECT  3.395 1.290 3.525 1.860 ;
        RECT  3.345 1.290 3.395 1.765 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.390 0.645 9.550 2.925 ;
        RECT  9.050 0.645 9.390 0.805 ;
        RECT  9.325 2.520 9.390 2.925 ;
        RECT  9.040 2.765 9.325 2.925 ;
        RECT  8.790 0.490 9.050 0.805 ;
        RECT  8.780 2.765 9.040 3.025 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.990 1.105 9.995 2.585 ;
        RECT  9.785 0.920 9.990 2.750 ;
        RECT  9.730 0.920 9.785 1.180 ;
        RECT  9.730 2.150 9.785 2.750 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.285 0.440 1.545 ;
        RECT  0.125 1.285 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.690 1.630 3.155 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.590 -0.250 10.120 0.250 ;
        RECT  9.330 -0.250 9.590 0.405 ;
        RECT  8.510 -0.250 9.330 0.250 ;
        RECT  8.250 -0.250 8.510 1.240 ;
        RECT  4.655 -0.250 8.250 0.250 ;
        RECT  4.055 -0.250 4.655 0.405 ;
        RECT  2.140 -0.250 4.055 0.250 ;
        RECT  1.880 -0.250 2.140 0.405 ;
        RECT  0.385 -0.250 1.880 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.590 3.440 10.120 3.940 ;
        RECT  9.330 3.285 9.590 3.940 ;
        RECT  8.530 3.440 9.330 3.940 ;
        RECT  8.370 2.380 8.530 3.940 ;
        RECT  8.230 2.380 8.370 2.640 ;
        RECT  6.425 3.440 8.370 3.940 ;
        RECT  6.165 3.115 6.425 3.940 ;
        RECT  4.705 3.440 6.165 3.940 ;
        RECT  3.765 3.055 4.705 3.940 ;
        RECT  2.205 3.440 3.765 3.940 ;
        RECT  1.945 3.285 2.205 3.940 ;
        RECT  0.535 3.440 1.945 3.940 ;
        RECT  0.275 2.500 0.535 3.940 ;
        RECT  0.000 3.440 0.275 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.080 1.105 9.205 2.120 ;
        RECT  9.045 1.105 9.080 2.345 ;
        RECT  8.820 1.105 9.045 1.365 ;
        RECT  8.820 1.960 9.045 2.345 ;
        RECT  7.715 1.960 8.820 2.120 ;
        RECT  8.065 1.560 8.670 1.720 ;
        RECT  7.905 1.280 8.065 1.720 ;
        RECT  7.870 0.770 7.970 1.030 ;
        RECT  7.655 2.405 7.915 2.665 ;
        RECT  6.825 1.280 7.905 1.440 ;
        RECT  7.710 0.470 7.870 1.030 ;
        RECT  7.455 1.910 7.715 2.170 ;
        RECT  5.245 0.470 7.710 0.630 ;
        RECT  7.540 2.505 7.655 2.665 ;
        RECT  7.380 2.505 7.540 2.935 ;
        RECT  5.230 2.775 7.380 2.935 ;
        RECT  7.030 0.810 7.290 1.095 ;
        RECT  7.005 1.620 7.165 2.595 ;
        RECT  6.365 0.810 7.030 0.970 ;
        RECT  6.905 1.620 7.005 1.880 ;
        RECT  5.575 2.435 7.005 2.595 ;
        RECT  6.725 1.150 6.825 1.440 ;
        RECT  6.725 2.095 6.825 2.255 ;
        RECT  6.565 1.150 6.725 2.255 ;
        RECT  6.205 0.810 6.365 2.060 ;
        RECT  5.585 0.810 6.205 0.970 ;
        RECT  5.925 1.150 6.025 1.310 ;
        RECT  5.925 2.095 6.025 2.255 ;
        RECT  5.765 1.150 5.925 2.255 ;
        RECT  4.565 1.465 5.765 1.625 ;
        RECT  5.425 0.810 5.585 1.285 ;
        RECT  5.415 2.160 5.575 2.595 ;
        RECT  4.905 1.125 5.425 1.285 ;
        RECT  4.845 2.160 5.415 2.320 ;
        RECT  5.085 0.470 5.245 0.945 ;
        RECT  5.070 2.515 5.230 2.935 ;
        RECT  4.225 1.805 5.080 1.965 ;
        RECT  4.745 0.585 4.905 1.285 ;
        RECT  4.685 2.160 4.845 2.860 ;
        RECT  3.845 0.585 4.745 0.745 ;
        RECT  3.405 2.700 4.685 2.860 ;
        RECT  4.405 0.925 4.565 1.625 ;
        RECT  3.505 0.925 4.405 1.085 ;
        RECT  4.125 1.265 4.225 2.415 ;
        RECT  4.065 1.265 4.125 2.465 ;
        RECT  3.965 1.265 4.065 1.425 ;
        RECT  3.865 2.205 4.065 2.465 ;
        RECT  3.685 0.470 3.845 0.745 ;
        RECT  2.785 0.470 3.685 0.630 ;
        RECT  3.345 0.845 3.505 1.085 ;
        RECT  3.245 2.170 3.405 2.910 ;
        RECT  2.825 0.845 3.345 1.005 ;
        RECT  2.455 2.170 3.245 2.330 ;
        RECT  3.065 3.100 3.245 3.260 ;
        RECT  3.005 1.185 3.165 1.445 ;
        RECT  2.905 2.510 3.065 3.260 ;
        RECT  2.455 1.285 3.005 1.445 ;
        RECT  1.395 2.510 2.905 2.670 ;
        RECT  2.665 0.845 2.825 1.085 ;
        RECT  2.525 0.445 2.785 0.630 ;
        RECT  2.565 2.850 2.725 3.110 ;
        RECT  2.095 0.925 2.665 1.085 ;
        RECT  1.620 2.850 2.565 3.010 ;
        RECT  2.485 0.470 2.525 0.630 ;
        RECT  2.325 0.470 2.485 0.745 ;
        RECT  2.295 1.285 2.455 2.330 ;
        RECT  0.955 0.585 2.325 0.745 ;
        RECT  2.285 1.645 2.295 2.330 ;
        RECT  1.715 1.645 2.285 1.805 ;
        RECT  1.935 0.925 2.095 1.425 ;
        RECT  1.835 1.165 1.935 1.425 ;
        RECT  1.555 1.645 1.715 1.910 ;
        RECT  1.360 2.850 1.620 3.045 ;
        RECT  1.375 0.975 1.395 1.135 ;
        RECT  1.375 2.270 1.395 2.670 ;
        RECT  1.215 0.975 1.375 2.670 ;
        RECT  0.935 2.850 1.360 3.010 ;
        RECT  1.135 0.975 1.215 1.135 ;
        RECT  1.185 2.270 1.215 2.670 ;
        RECT  1.135 2.270 1.185 2.530 ;
        RECT  0.955 1.335 1.035 1.595 ;
        RECT  0.935 0.585 0.955 1.595 ;
        RECT  0.795 0.585 0.935 3.010 ;
        RECT  0.775 1.335 0.795 3.010 ;
    END
END DFFNSRX1

MACRO DFFNSRXL
    CLASS CORE ;
    FOREIGN DFFNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.725 2.890 8.185 3.260 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.700 3.885 1.960 ;
        RECT  3.530 1.290 3.555 1.960 ;
        RECT  3.395 1.290 3.530 1.860 ;
        RECT  3.345 1.290 3.395 1.765 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.390 0.645 9.550 2.970 ;
        RECT  9.055 0.645 9.390 0.805 ;
        RECT  9.325 2.520 9.390 2.970 ;
        RECT  9.070 2.810 9.325 2.970 ;
        RECT  8.810 2.810 9.070 3.100 ;
        RECT  8.795 0.545 9.055 0.805 ;
        END
        ANTENNADIFFAREA     0.2135 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.990 0.920 9.995 2.585 ;
        RECT  9.785 0.920 9.990 2.880 ;
        RECT  9.735 0.920 9.785 1.180 ;
        RECT  9.730 2.620 9.785 2.880 ;
        END
        ANTENNADIFFAREA     0.2135 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.285 0.440 1.545 ;
        RECT  0.125 1.285 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.690 1.645 3.165 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.565 -0.250 10.120 0.250 ;
        RECT  9.305 -0.250 9.565 0.405 ;
        RECT  8.485 -0.250 9.305 0.250 ;
        RECT  8.225 -0.250 8.485 1.240 ;
        RECT  4.645 -0.250 8.225 0.250 ;
        RECT  4.045 -0.250 4.645 0.405 ;
        RECT  2.140 -0.250 4.045 0.250 ;
        RECT  1.880 -0.250 2.140 0.405 ;
        RECT  0.385 -0.250 1.880 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.590 3.440 10.120 3.940 ;
        RECT  9.330 3.285 9.590 3.940 ;
        RECT  8.530 3.440 9.330 3.940 ;
        RECT  8.370 2.460 8.530 3.940 ;
        RECT  8.260 2.460 8.370 2.720 ;
        RECT  6.425 3.440 8.370 3.940 ;
        RECT  6.165 3.115 6.425 3.940 ;
        RECT  4.705 3.440 6.165 3.940 ;
        RECT  3.765 3.055 4.705 3.940 ;
        RECT  2.205 3.440 3.765 3.940 ;
        RECT  1.945 3.285 2.205 3.940 ;
        RECT  0.505 3.440 1.945 3.940 ;
        RECT  0.245 2.500 0.505 3.940 ;
        RECT  0.000 3.440 0.245 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.100 1.095 9.180 2.120 ;
        RECT  9.020 1.095 9.100 2.355 ;
        RECT  8.795 1.095 9.020 1.355 ;
        RECT  8.840 1.960 9.020 2.355 ;
        RECT  7.455 1.960 8.840 2.120 ;
        RECT  8.410 1.510 8.670 1.770 ;
        RECT  7.895 1.510 8.410 1.670 ;
        RECT  7.845 0.845 7.945 1.105 ;
        RECT  7.655 2.405 7.915 2.665 ;
        RECT  7.735 1.365 7.895 1.670 ;
        RECT  7.685 0.470 7.845 1.105 ;
        RECT  6.825 1.365 7.735 1.525 ;
        RECT  5.245 0.470 7.685 0.630 ;
        RECT  7.540 2.505 7.655 2.665 ;
        RECT  7.380 2.505 7.540 2.935 ;
        RECT  5.230 2.775 7.380 2.935 ;
        RECT  7.005 0.810 7.265 1.095 ;
        RECT  7.010 1.720 7.170 2.595 ;
        RECT  6.905 1.720 7.010 1.880 ;
        RECT  5.575 2.435 7.010 2.595 ;
        RECT  6.365 0.810 7.005 0.970 ;
        RECT  6.725 1.150 6.825 1.525 ;
        RECT  6.725 2.095 6.825 2.255 ;
        RECT  6.565 1.150 6.725 2.255 ;
        RECT  6.205 0.810 6.365 2.060 ;
        RECT  5.585 0.810 6.205 0.970 ;
        RECT  5.925 1.150 6.025 1.310 ;
        RECT  5.925 2.095 6.025 2.255 ;
        RECT  5.765 1.150 5.925 2.255 ;
        RECT  4.565 1.465 5.765 1.625 ;
        RECT  5.425 0.810 5.585 1.285 ;
        RECT  5.415 2.160 5.575 2.595 ;
        RECT  4.905 1.125 5.425 1.285 ;
        RECT  4.890 2.160 5.415 2.320 ;
        RECT  5.085 0.470 5.245 0.945 ;
        RECT  5.070 2.515 5.230 2.935 ;
        RECT  4.225 1.805 5.070 1.965 ;
        RECT  4.745 0.585 4.905 1.285 ;
        RECT  4.730 2.160 4.890 2.755 ;
        RECT  3.845 0.585 4.745 0.745 ;
        RECT  3.405 2.595 4.730 2.755 ;
        RECT  4.405 0.925 4.565 1.625 ;
        RECT  3.505 0.925 4.405 1.085 ;
        RECT  4.065 1.265 4.225 2.415 ;
        RECT  3.955 1.265 4.065 1.425 ;
        RECT  3.865 2.255 4.065 2.415 ;
        RECT  3.685 0.470 3.845 0.745 ;
        RECT  2.785 0.470 3.685 0.630 ;
        RECT  3.345 0.845 3.505 1.085 ;
        RECT  3.245 2.170 3.405 2.910 ;
        RECT  2.825 0.845 3.345 1.005 ;
        RECT  2.445 2.170 3.245 2.330 ;
        RECT  3.065 3.100 3.245 3.260 ;
        RECT  3.005 1.185 3.165 1.445 ;
        RECT  2.905 2.510 3.065 3.260 ;
        RECT  2.445 1.285 3.005 1.445 ;
        RECT  1.375 2.510 2.905 2.670 ;
        RECT  2.665 0.845 2.825 1.085 ;
        RECT  2.525 0.445 2.785 0.630 ;
        RECT  2.565 2.850 2.725 3.110 ;
        RECT  2.045 0.925 2.665 1.085 ;
        RECT  1.625 2.850 2.565 3.010 ;
        RECT  2.485 0.470 2.525 0.630 ;
        RECT  2.325 0.470 2.485 0.745 ;
        RECT  2.285 1.285 2.445 2.330 ;
        RECT  0.945 0.585 2.325 0.745 ;
        RECT  1.685 1.645 2.285 1.805 ;
        RECT  1.885 0.925 2.045 1.425 ;
        RECT  1.525 1.645 1.685 1.910 ;
        RECT  1.415 2.850 1.625 3.045 ;
        RECT  1.365 2.865 1.415 3.045 ;
        RECT  1.345 0.925 1.395 1.185 ;
        RECT  1.345 2.270 1.375 2.670 ;
        RECT  0.985 2.865 1.365 3.025 ;
        RECT  1.185 0.925 1.345 2.670 ;
        RECT  1.135 0.925 1.185 1.185 ;
        RECT  0.945 1.335 0.985 3.025 ;
        RECT  0.825 0.585 0.945 3.025 ;
        RECT  0.785 0.585 0.825 1.545 ;
    END
END DFFNSRXL

MACRO DFFSRX4
    CLASS CORE ;
    FOREIGN DFFSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.640 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.145 2.930 12.295 3.220 ;
        RECT  11.935 2.520 12.145 3.220 ;
        RECT  11.860 2.520 11.935 2.810 ;
        END
        ANTENNAGATEAREA     0.3250 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.285 2.110 4.475 2.400 ;
        RECT  4.265 1.620 4.285 2.400 ;
        RECT  4.125 1.620 4.265 2.270 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.455 0.595 14.615 2.320 ;
        RECT  12.955 0.595 14.455 0.755 ;
        RECT  13.670 2.160 14.455 2.320 ;
        RECT  13.670 2.520 13.675 3.220 ;
        RECT  13.465 2.160 13.670 3.220 ;
        RECT  13.400 2.160 13.465 3.100 ;
        RECT  12.695 0.595 12.955 1.195 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.320 1.290 15.515 1.990 ;
        RECT  15.305 1.085 15.320 1.990 ;
        RECT  14.955 1.085 15.305 2.745 ;
        RECT  14.845 0.645 14.955 2.745 ;
        RECT  14.795 0.645 14.845 1.245 ;
        RECT  14.680 2.505 14.845 2.745 ;
        RECT  14.420 2.505 14.680 3.105 ;
        RECT  14.385 2.745 14.420 2.995 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.335 2.025 ;
        END
        ANTENNAGATEAREA     0.2457 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.635 3.505 1.895 ;
        RECT  2.635 1.700 3.345 1.860 ;
        RECT  2.425 1.700 2.635 1.990 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.515 -0.250 15.640 0.250 ;
        RECT  15.255 -0.250 15.515 0.795 ;
        RECT  14.455 -0.250 15.255 0.250 ;
        RECT  14.195 -0.250 14.455 0.405 ;
        RECT  13.505 -0.250 14.195 0.250 ;
        RECT  13.245 -0.250 13.505 0.405 ;
        RECT  12.445 -0.250 13.245 0.250 ;
        RECT  12.185 -0.250 12.445 1.165 ;
        RECT  11.385 -0.250 12.185 0.250 ;
        RECT  11.125 -0.250 11.385 1.135 ;
        RECT  3.945 -0.250 11.125 0.250 ;
        RECT  3.685 -0.250 3.945 0.405 ;
        RECT  2.450 -0.250 3.685 0.250 ;
        RECT  2.190 -0.250 2.450 0.405 ;
        RECT  0.525 -0.250 2.190 0.250 ;
        RECT  0.265 -0.250 0.525 0.905 ;
        RECT  0.000 -0.250 0.265 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.205 3.440 15.640 3.940 ;
        RECT  14.945 2.955 15.205 3.940 ;
        RECT  14.170 3.440 14.945 3.940 ;
        RECT  13.910 2.600 14.170 3.940 ;
        RECT  13.140 3.440 13.910 3.940 ;
        RECT  12.880 2.445 13.140 3.940 ;
        RECT  9.880 3.440 12.880 3.940 ;
        RECT  9.280 3.285 9.880 3.940 ;
        RECT  6.600 3.440 9.280 3.940 ;
        RECT  6.340 3.105 6.600 3.940 ;
        RECT  5.010 3.440 6.340 3.940 ;
        RECT  4.410 3.105 5.010 3.940 ;
        RECT  2.570 3.440 4.410 3.940 ;
        RECT  2.310 3.115 2.570 3.940 ;
        RECT  0.435 3.440 2.310 3.940 ;
        RECT  0.175 2.610 0.435 3.940 ;
        RECT  0.000 3.440 0.175 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.100 0.955 14.260 1.980 ;
        RECT  13.645 0.955 14.100 1.115 ;
        RECT  12.620 1.820 14.100 1.980 ;
        RECT  12.280 1.470 13.805 1.630 ;
        RECT  12.460 1.820 12.620 2.735 ;
        RECT  12.360 2.080 12.460 2.735 ;
        RECT  11.460 2.080 12.360 2.240 ;
        RECT  12.115 1.470 12.280 1.900 ;
        RECT  10.475 1.740 12.115 1.900 ;
        RECT  11.835 0.495 11.935 1.435 ;
        RECT  11.675 0.495 11.835 1.560 ;
        RECT  11.630 2.810 11.680 3.070 ;
        RECT  10.815 1.400 11.675 1.560 ;
        RECT  11.420 2.810 11.630 3.205 ;
        RECT  11.200 2.080 11.460 2.340 ;
        RECT  10.460 3.045 11.420 3.205 ;
        RECT  10.950 2.570 10.955 2.765 ;
        RECT  10.790 2.520 10.950 2.780 ;
        RECT  10.655 0.475 10.815 1.560 ;
        RECT  7.555 2.605 10.790 2.765 ;
        RECT  10.540 0.475 10.655 0.635 ;
        RECT  10.475 2.265 10.610 2.425 ;
        RECT  10.280 0.470 10.540 0.635 ;
        RECT  10.315 0.815 10.475 2.425 ;
        RECT  10.300 2.945 10.460 3.205 ;
        RECT  8.835 0.815 10.315 0.975 ;
        RECT  8.510 2.265 10.315 2.425 ;
        RECT  7.150 2.945 10.300 3.105 ;
        RECT  8.160 0.475 10.280 0.635 ;
        RECT  9.975 1.160 10.135 2.065 ;
        RECT  8.345 1.160 9.975 1.320 ;
        RECT  7.730 1.905 9.975 2.065 ;
        RECT  9.530 1.535 9.790 1.725 ;
        RECT  7.030 1.535 9.530 1.695 ;
        RECT  8.250 2.245 8.510 2.425 ;
        RECT  7.795 1.025 8.345 1.320 ;
        RECT  7.900 0.475 8.160 0.735 ;
        RECT  7.070 0.525 7.900 0.685 ;
        RECT  7.405 1.025 7.795 1.285 ;
        RECT  7.570 1.905 7.730 2.245 ;
        RECT  5.240 2.085 7.570 2.245 ;
        RECT  7.395 2.425 7.555 2.765 ;
        RECT  6.495 1.025 7.405 1.185 ;
        RECT  5.405 2.425 7.395 2.585 ;
        RECT  6.990 2.765 7.150 3.105 ;
        RECT  6.810 0.495 7.070 0.755 ;
        RECT  6.870 1.370 7.030 1.695 ;
        RECT  6.890 2.765 6.990 2.940 ;
        RECT  6.050 2.765 6.890 2.925 ;
        RECT  4.985 1.370 6.870 1.530 ;
        RECT  6.235 0.925 6.495 1.185 ;
        RECT  6.130 1.715 6.390 1.890 ;
        RECT  5.530 1.025 6.235 1.185 ;
        RECT  4.870 1.730 6.130 1.890 ;
        RECT  5.780 2.765 6.050 2.940 ;
        RECT  5.430 0.885 5.530 1.185 ;
        RECT  5.270 0.595 5.430 1.185 ;
        RECT  5.245 2.425 5.405 2.875 ;
        RECT  3.445 0.595 5.270 0.755 ;
        RECT  3.260 2.715 5.245 2.875 ;
        RECT  4.825 0.935 4.985 1.530 ;
        RECT  4.870 2.355 4.980 2.515 ;
        RECT  4.710 1.730 4.870 2.515 ;
        RECT  3.940 0.935 4.825 1.095 ;
        RECT  4.635 1.730 4.710 1.910 ;
        RECT  4.475 1.275 4.635 1.910 ;
        RECT  4.245 1.275 4.475 1.435 ;
        RECT  3.850 0.935 3.940 1.435 ;
        RECT  3.780 0.935 3.850 2.535 ;
        RECT  3.690 1.275 3.780 2.535 ;
        RECT  2.915 3.060 3.725 3.220 ;
        RECT  3.115 1.275 3.690 1.435 ;
        RECT  3.560 2.085 3.690 2.535 ;
        RECT  2.815 2.085 3.560 2.245 ;
        RECT  3.285 0.595 3.445 1.090 ;
        RECT  2.565 0.930 3.285 1.090 ;
        RECT  3.100 2.425 3.260 2.875 ;
        RECT  1.975 0.585 3.100 0.745 ;
        RECT  1.975 2.425 3.100 2.585 ;
        RECT  2.755 2.770 2.915 3.220 ;
        RECT  1.620 2.770 2.755 2.930 ;
        RECT  2.405 0.930 2.565 1.505 ;
        RECT  2.305 1.245 2.405 1.505 ;
        RECT  1.975 1.345 2.025 1.605 ;
        RECT  1.815 0.585 1.975 2.585 ;
        RECT  1.765 1.345 1.815 1.940 ;
        RECT  1.035 1.780 1.765 1.940 ;
        RECT  1.020 2.240 1.620 2.930 ;
        RECT  1.325 0.555 1.425 1.155 ;
        RECT  1.165 0.555 1.325 1.485 ;
        RECT  0.685 1.325 1.165 1.485 ;
        RECT  0.875 1.730 1.035 1.990 ;
        RECT  0.685 2.240 1.020 2.400 ;
        RECT  0.525 1.325 0.685 2.400 ;
    END
END DFFSRX4

MACRO DFFSRX2
    CLASS CORE ;
    FOREIGN DFFSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.795 2.925 8.355 3.225 ;
        END
        ANTENNAGATEAREA     0.1859 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.615 1.610 4.015 2.035 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.765 1.115 10.925 2.060 ;
        RECT  10.340 1.115 10.765 1.275 ;
        RECT  10.340 1.900 10.765 2.060 ;
        RECT  10.080 0.675 10.340 1.275 ;
        RECT  10.180 1.900 10.340 3.220 ;
        RECT  10.080 2.255 10.180 3.220 ;
        RECT  9.785 2.930 10.080 3.220 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.370 0.695 11.375 2.585 ;
        RECT  11.110 0.695 11.370 2.895 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.850 0.445 2.480 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.715 1.645 3.095 1.990 ;
        END
        ANTENNAGATEAREA     0.0637 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.855 -0.250 11.500 0.250 ;
        RECT  10.595 -0.250 10.855 0.865 ;
        RECT  9.715 -0.250 10.595 0.250 ;
        RECT  8.775 -0.250 9.715 0.405 ;
        RECT  3.160 -0.250 8.775 0.250 ;
        RECT  2.900 -0.250 3.160 0.405 ;
        RECT  2.015 -0.250 2.900 0.250 ;
        RECT  1.755 -0.250 2.015 0.405 ;
        RECT  0.385 -0.250 1.755 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.860 3.440 11.500 3.940 ;
        RECT  10.600 2.255 10.860 3.940 ;
        RECT  9.605 3.440 10.600 3.940 ;
        RECT  9.345 2.825 9.605 3.940 ;
        RECT  6.165 3.440 9.345 3.940 ;
        RECT  5.905 3.285 6.165 3.940 ;
        RECT  4.405 3.440 5.905 3.940 ;
        RECT  3.465 3.055 4.405 3.940 ;
        RECT  2.030 3.440 3.465 3.940 ;
        RECT  1.770 2.900 2.030 3.940 ;
        RECT  0.390 3.440 1.770 3.940 ;
        RECT  0.130 2.810 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.610 1.455 10.585 1.715 ;
        RECT  9.450 1.135 9.610 2.615 ;
        RECT  9.360 1.135 9.450 1.295 ;
        RECT  9.065 2.455 9.450 2.615 ;
        RECT  9.100 1.035 9.360 1.295 ;
        RECT  9.170 1.545 9.265 1.805 ;
        RECT  9.010 1.545 9.170 2.190 ;
        RECT  8.805 2.455 9.065 2.730 ;
        RECT  9.005 1.545 9.010 1.805 ;
        RECT  7.360 2.030 9.010 2.190 ;
        RECT  8.185 2.455 8.805 2.615 ;
        RECT  8.190 0.475 8.450 0.755 ;
        RECT  5.660 0.475 8.190 0.635 ;
        RECT  7.925 2.405 8.185 2.665 ;
        RECT  7.805 0.815 7.965 1.795 ;
        RECT  6.600 0.815 7.805 0.975 ;
        RECT  7.615 1.635 7.805 1.795 ;
        RECT  7.465 1.155 7.625 1.415 ;
        RECT  7.350 2.785 7.610 3.105 ;
        RECT  7.360 1.250 7.465 1.415 ;
        RECT  7.200 1.250 7.360 2.190 ;
        RECT  4.875 2.945 7.350 3.105 ;
        RECT  7.115 1.250 7.200 1.920 ;
        RECT  6.305 1.760 7.115 1.920 ;
        RECT  6.825 2.265 6.925 2.525 ;
        RECT  6.665 2.265 6.825 2.765 ;
        RECT  4.530 2.605 6.665 2.765 ;
        RECT  6.450 0.815 6.600 1.505 ;
        RECT  6.440 0.815 6.450 1.580 ;
        RECT  6.190 1.320 6.440 1.580 ;
        RECT  6.145 1.760 6.305 2.360 ;
        RECT  5.965 1.420 6.190 1.580 ;
        RECT  6.010 0.855 6.170 1.015 ;
        RECT  5.845 0.855 6.010 1.240 ;
        RECT  5.805 1.420 5.965 2.325 ;
        RECT  5.625 1.080 5.845 1.240 ;
        RECT  4.795 2.165 5.805 2.325 ;
        RECT  5.500 0.475 5.660 0.900 ;
        RECT  5.465 1.080 5.625 1.985 ;
        RECT  5.400 0.740 5.500 0.900 ;
        RECT  5.100 1.080 5.465 1.240 ;
        RECT  4.940 0.475 5.100 1.240 ;
        RECT  3.500 0.475 4.940 0.635 ;
        RECT  4.730 1.420 4.795 2.325 ;
        RECT  4.635 0.815 4.730 2.325 ;
        RECT  4.570 0.815 4.635 1.580 ;
        RECT  3.840 0.815 4.570 0.975 ;
        RECT  4.370 2.605 4.530 2.870 ;
        RECT  4.355 1.760 4.455 1.920 ;
        RECT  2.715 2.710 4.370 2.870 ;
        RECT  4.195 1.155 4.355 2.375 ;
        RECT  4.020 1.155 4.195 1.315 ;
        RECT  4.190 2.215 4.195 2.375 ;
        RECT  3.930 2.215 4.190 2.475 ;
        RECT  3.680 0.815 3.840 1.430 ;
        RECT  3.435 1.270 3.680 1.430 ;
        RECT  3.340 0.475 3.500 1.090 ;
        RECT  3.275 1.270 3.435 2.355 ;
        RECT  1.955 0.930 3.340 1.090 ;
        RECT  2.360 1.270 3.275 1.430 ;
        RECT  2.915 2.195 3.275 2.355 ;
        RECT  2.985 3.050 3.245 3.240 ;
        RECT  2.370 3.050 2.985 3.210 ;
        RECT  2.555 2.215 2.715 2.870 ;
        RECT  2.390 0.490 2.650 0.750 ;
        RECT  1.825 2.215 2.555 2.375 ;
        RECT  1.425 0.590 2.390 0.750 ;
        RECT  2.210 2.560 2.370 3.210 ;
        RECT  2.200 1.270 2.360 2.035 ;
        RECT  1.310 2.560 2.210 2.720 ;
        RECT  1.795 0.930 1.955 1.365 ;
        RECT  1.665 2.025 1.825 2.375 ;
        RECT  1.695 1.105 1.795 1.365 ;
        RECT  1.425 2.025 1.665 2.185 ;
        RECT  1.265 0.590 1.425 2.185 ;
        RECT  1.000 2.440 1.310 2.720 ;
        RECT  0.970 1.925 1.265 2.185 ;
        RECT  0.885 0.825 1.045 1.085 ;
        RECT  0.790 2.440 1.000 2.600 ;
        RECT  0.790 0.925 0.885 1.085 ;
        RECT  0.630 0.925 0.790 2.600 ;
    END
END DFFSRX2

MACRO DFFSRX1
    CLASS CORE ;
    FOREIGN DFFSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.050 2.520 8.155 2.810 ;
        RECT  7.890 2.520 8.050 3.175 ;
        RECT  7.790 2.915 7.890 3.175 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.765 4.075 2.065 ;
        RECT  3.715 1.700 4.015 2.065 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.530 2.335 9.535 2.810 ;
        RECT  9.370 0.645 9.530 2.810 ;
        RECT  9.325 0.645 9.370 0.945 ;
        RECT  9.325 2.335 9.370 2.810 ;
        RECT  9.065 0.645 9.325 0.805 ;
        RECT  9.080 2.595 9.325 2.810 ;
        RECT  8.820 2.595 9.080 3.195 ;
        RECT  8.805 0.545 9.065 0.805 ;
        END
        ANTENNADIFFAREA     0.3838 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.990 0.920 9.995 2.585 ;
        RECT  9.785 0.920 9.990 2.750 ;
        RECT  9.735 0.920 9.785 1.180 ;
        RECT  9.730 2.150 9.785 2.750 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 1.990 0.455 2.250 ;
        RECT  0.195 1.700 0.405 2.250 ;
        RECT  0.125 1.700 0.195 1.990 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.625 1.695 3.095 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.595 -0.250 10.120 0.250 ;
        RECT  9.335 -0.250 9.595 0.405 ;
        RECT  8.515 -0.250 9.335 0.250 ;
        RECT  8.255 -0.250 8.515 0.405 ;
        RECT  3.760 -0.250 8.255 0.250 ;
        RECT  3.500 -0.250 3.760 0.405 ;
        RECT  2.065 -0.250 3.500 0.250 ;
        RECT  1.805 -0.250 2.065 0.405 ;
        RECT  0.395 -0.250 1.805 0.250 ;
        RECT  0.135 -0.250 0.395 0.405 ;
        RECT  0.000 -0.250 0.135 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.590 3.440 10.120 3.940 ;
        RECT  9.330 3.285 9.590 3.940 ;
        RECT  8.510 3.440 9.330 3.940 ;
        RECT  8.250 3.285 8.510 3.940 ;
        RECT  6.245 3.440 8.250 3.940 ;
        RECT  5.985 3.285 6.245 3.940 ;
        RECT  4.390 3.440 5.985 3.940 ;
        RECT  3.450 2.975 4.390 3.940 ;
        RECT  2.000 3.440 3.450 3.940 ;
        RECT  1.840 2.900 2.000 3.940 ;
        RECT  0.385 3.440 1.840 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.100 1.635 9.190 1.895 ;
        RECT  9.080 1.120 9.100 2.085 ;
        RECT  8.940 1.120 9.080 2.345 ;
        RECT  8.825 1.120 8.940 1.380 ;
        RECT  8.820 1.910 8.940 2.345 ;
        RECT  7.740 1.910 8.820 2.070 ;
        RECT  8.570 1.560 8.760 1.720 ;
        RECT  8.410 1.275 8.570 1.720 ;
        RECT  7.040 1.275 8.410 1.435 ;
        RECT  8.010 0.805 8.110 1.065 ;
        RECT  7.850 0.475 8.010 1.065 ;
        RECT  5.440 0.475 7.850 0.635 ;
        RECT  7.480 1.825 7.740 2.085 ;
        RECT  7.515 2.285 7.615 2.545 ;
        RECT  7.355 2.285 7.515 3.100 ;
        RECT  7.220 0.815 7.380 1.095 ;
        RECT  5.150 2.940 7.355 3.100 ;
        RECT  6.290 0.815 7.220 0.975 ;
        RECT  6.970 1.615 7.070 1.775 ;
        RECT  6.755 1.175 7.040 1.435 ;
        RECT  6.810 1.615 6.970 2.755 ;
        RECT  4.760 2.595 6.810 2.755 ;
        RECT  6.630 1.275 6.755 1.435 ;
        RECT  6.470 1.275 6.630 2.385 ;
        RECT  6.030 2.125 6.470 2.385 ;
        RECT  6.130 0.815 6.290 1.920 ;
        RECT  5.900 1.660 6.130 1.920 ;
        RECT  5.790 0.815 5.950 1.285 ;
        RECT  5.840 1.760 5.900 1.920 ;
        RECT  5.680 1.760 5.840 2.415 ;
        RECT  5.480 1.125 5.790 1.285 ;
        RECT  5.120 2.255 5.680 2.415 ;
        RECT  5.320 1.125 5.480 2.050 ;
        RECT  5.280 0.475 5.440 0.945 ;
        RECT  5.100 1.125 5.320 1.285 ;
        RECT  4.990 2.940 5.150 3.225 ;
        RECT  4.960 1.465 5.120 2.415 ;
        RECT  4.940 0.590 5.100 1.285 ;
        RECT  4.830 2.965 4.990 3.225 ;
        RECT  4.760 1.465 4.960 1.625 ;
        RECT  3.095 0.590 4.940 0.750 ;
        RECT  4.600 0.930 4.760 1.625 ;
        RECT  4.425 1.850 4.760 2.110 ;
        RECT  4.600 2.595 4.760 2.775 ;
        RECT  3.470 0.930 4.600 1.090 ;
        RECT  2.830 2.615 4.600 2.775 ;
        RECT  4.420 1.850 4.425 2.425 ;
        RECT  4.260 1.270 4.420 2.425 ;
        RECT  4.040 1.270 4.260 1.430 ;
        RECT  3.880 2.265 4.260 2.425 ;
        RECT  3.310 0.930 3.470 2.355 ;
        RECT  2.410 1.270 3.310 1.430 ;
        RECT  2.865 2.195 3.310 2.355 ;
        RECT  2.985 3.050 3.245 3.260 ;
        RECT  2.935 0.590 3.095 1.090 ;
        RECT  2.345 3.050 2.985 3.210 ;
        RECT  1.925 0.930 2.935 1.090 ;
        RECT  2.685 2.615 2.830 2.870 ;
        RECT  2.525 2.215 2.685 2.870 ;
        RECT  1.430 0.590 2.660 0.750 ;
        RECT  1.695 2.215 2.525 2.375 ;
        RECT  2.250 1.270 2.410 2.035 ;
        RECT  2.185 2.560 2.345 3.210 ;
        RECT  2.150 1.775 2.250 2.035 ;
        RECT  1.320 2.560 2.185 2.720 ;
        RECT  1.765 0.930 1.925 1.455 ;
        RECT  1.665 1.195 1.765 1.455 ;
        RECT  1.535 2.160 1.695 2.375 ;
        RECT  1.345 2.160 1.535 2.320 ;
        RECT  1.345 0.590 1.430 1.475 ;
        RECT  1.270 0.590 1.345 2.320 ;
        RECT  1.055 2.500 1.320 2.720 ;
        RECT  1.145 1.265 1.270 2.320 ;
        RECT  1.085 1.265 1.145 1.525 ;
        RECT  1.050 2.060 1.145 2.320 ;
        RECT  0.925 0.820 1.085 1.080 ;
        RECT  0.870 2.500 1.055 2.660 ;
        RECT  0.870 0.920 0.925 1.080 ;
        RECT  0.710 0.920 0.870 2.660 ;
    END
END DFFSRX1

MACRO DFFSRXL
    CLASS CORE ;
    FOREIGN DFFSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.010 2.520 8.155 2.810 ;
        RECT  7.850 2.520 8.010 3.175 ;
        RECT  7.750 2.915 7.850 3.175 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 1.700 4.015 1.990 ;
        RECT  3.615 1.700 3.970 2.065 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.515 1.105 9.535 1.355 ;
        RECT  9.515 2.335 9.535 2.810 ;
        RECT  9.355 0.645 9.515 2.810 ;
        RECT  9.325 0.645 9.355 1.355 ;
        RECT  9.325 2.335 9.355 2.810 ;
        RECT  9.055 0.645 9.325 0.805 ;
        RECT  9.040 2.650 9.325 2.810 ;
        RECT  8.795 0.545 9.055 0.805 ;
        RECT  8.830 2.650 9.040 3.025 ;
        RECT  8.780 2.765 8.830 3.025 ;
        END
        ANTENNADIFFAREA     0.2231 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.985 0.920 9.995 2.400 ;
        RECT  9.735 0.920 9.985 2.580 ;
        RECT  9.725 2.320 9.735 2.580 ;
        END
        ANTENNADIFFAREA     0.2199 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.365 1.990 0.415 2.250 ;
        RECT  0.155 1.700 0.365 2.250 ;
        RECT  0.125 1.700 0.155 2.175 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.625 1.695 3.095 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.565 -0.250 10.120 0.250 ;
        RECT  9.305 -0.250 9.565 0.405 ;
        RECT  8.460 -0.250 9.305 0.250 ;
        RECT  8.200 -0.250 8.460 0.405 ;
        RECT  3.720 -0.250 8.200 0.250 ;
        RECT  3.460 -0.250 3.720 0.405 ;
        RECT  2.125 -0.250 3.460 0.250 ;
        RECT  1.865 -0.250 2.125 0.405 ;
        RECT  0.385 -0.250 1.865 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.565 3.440 10.120 3.940 ;
        RECT  9.305 3.285 9.565 3.940 ;
        RECT  8.470 3.440 9.305 3.940 ;
        RECT  8.210 3.285 8.470 3.940 ;
        RECT  6.205 3.440 8.210 3.940 ;
        RECT  5.945 3.285 6.205 3.940 ;
        RECT  4.350 3.440 5.945 3.940 ;
        RECT  3.410 3.055 4.350 3.940 ;
        RECT  1.960 3.440 3.410 3.940 ;
        RECT  1.800 2.900 1.960 3.940 ;
        RECT  0.385 3.440 1.800 3.940 ;
        RECT  0.125 2.840 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.060 1.635 9.150 1.895 ;
        RECT  9.040 1.120 9.060 2.085 ;
        RECT  8.900 1.120 9.040 2.345 ;
        RECT  8.795 1.120 8.900 1.380 ;
        RECT  8.780 1.910 8.900 2.345 ;
        RECT  7.700 1.910 8.780 2.070 ;
        RECT  8.530 1.560 8.720 1.720 ;
        RECT  8.370 1.275 8.530 1.720 ;
        RECT  7.000 1.275 8.370 1.435 ;
        RECT  7.970 0.805 8.070 1.065 ;
        RECT  7.810 0.475 7.970 1.065 ;
        RECT  5.400 0.475 7.810 0.635 ;
        RECT  7.440 1.825 7.700 2.085 ;
        RECT  7.475 2.285 7.575 2.545 ;
        RECT  7.315 2.285 7.475 3.100 ;
        RECT  7.180 0.815 7.340 1.095 ;
        RECT  5.110 2.940 7.315 3.100 ;
        RECT  6.305 0.815 7.180 0.975 ;
        RECT  6.990 1.615 7.095 1.775 ;
        RECT  6.715 1.175 7.000 1.435 ;
        RECT  6.830 1.615 6.990 2.755 ;
        RECT  4.720 2.595 6.830 2.755 ;
        RECT  6.645 1.275 6.715 1.435 ;
        RECT  6.485 1.275 6.645 2.390 ;
        RECT  5.990 2.130 6.485 2.390 ;
        RECT  6.145 0.815 6.305 1.870 ;
        RECT  5.800 1.710 6.145 1.870 ;
        RECT  5.910 0.865 5.960 1.025 ;
        RECT  5.700 0.865 5.910 1.420 ;
        RECT  5.640 1.710 5.800 2.415 ;
        RECT  5.440 1.260 5.700 1.420 ;
        RECT  5.065 2.255 5.640 2.415 ;
        RECT  5.280 1.260 5.440 2.050 ;
        RECT  5.240 0.475 5.400 1.075 ;
        RECT  5.060 1.260 5.280 1.420 ;
        RECT  4.950 2.940 5.110 3.210 ;
        RECT  4.905 1.615 5.065 2.415 ;
        RECT  4.900 0.590 5.060 1.420 ;
        RECT  4.785 3.050 4.950 3.210 ;
        RECT  4.720 1.615 4.905 1.775 ;
        RECT  3.035 0.590 4.900 0.750 ;
        RECT  4.385 2.005 4.725 2.165 ;
        RECT  4.560 0.930 4.720 1.775 ;
        RECT  4.560 2.595 4.720 2.870 ;
        RECT  3.435 0.930 4.560 1.090 ;
        RECT  2.645 2.710 4.560 2.870 ;
        RECT  4.380 2.005 4.385 2.425 ;
        RECT  4.220 1.270 4.380 2.425 ;
        RECT  3.890 1.270 4.220 1.430 ;
        RECT  3.840 2.265 4.220 2.425 ;
        RECT  3.275 0.930 3.435 2.355 ;
        RECT  2.370 1.270 3.275 1.430 ;
        RECT  2.825 2.195 3.275 2.355 ;
        RECT  3.155 3.100 3.205 3.260 ;
        RECT  2.945 3.050 3.155 3.260 ;
        RECT  2.875 0.590 3.035 1.090 ;
        RECT  2.305 3.050 2.945 3.210 ;
        RECT  1.915 0.930 2.875 1.090 ;
        RECT  1.460 0.590 2.650 0.750 ;
        RECT  2.485 2.215 2.645 2.870 ;
        RECT  1.755 2.215 2.485 2.375 ;
        RECT  2.210 1.270 2.370 2.035 ;
        RECT  2.145 2.560 2.305 3.210 ;
        RECT  2.110 1.775 2.210 2.035 ;
        RECT  1.280 2.560 2.145 2.720 ;
        RECT  1.755 0.930 1.915 1.455 ;
        RECT  1.655 1.195 1.755 1.455 ;
        RECT  1.595 2.100 1.755 2.375 ;
        RECT  1.220 2.100 1.595 2.260 ;
        RECT  1.300 0.590 1.460 1.420 ;
        RECT  1.220 1.260 1.300 1.420 ;
        RECT  1.015 2.485 1.280 2.720 ;
        RECT  1.050 1.260 1.220 2.260 ;
        RECT  0.915 0.820 1.075 1.080 ;
        RECT  0.960 2.000 1.050 2.260 ;
        RECT  0.775 2.485 1.015 2.645 ;
        RECT  0.775 0.920 0.915 1.080 ;
        RECT  0.615 0.920 0.775 2.645 ;
    END
END DFFSRXL

MACRO DFFSX4
    CLASS CORE ;
    FOREIGN DFFSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.695 1.430 7.780 1.690 ;
        RECT  7.525 1.430 7.695 1.990 ;
        RECT  7.365 1.430 7.525 3.260 ;
        RECT  6.865 3.100 7.365 3.260 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.725 1.375 10.885 2.350 ;
        RECT  10.425 1.375 10.725 1.535 ;
        RECT  10.285 2.190 10.725 2.350 ;
        RECT  10.265 0.585 10.425 1.535 ;
        RECT  10.125 2.190 10.285 3.105 ;
        RECT  9.190 0.585 10.265 0.745 ;
        RECT  8.735 2.945 10.125 3.105 ;
        RECT  8.930 0.535 9.190 1.135 ;
        RECT  8.865 0.695 8.930 0.945 ;
        RECT  8.615 2.605 8.735 3.205 ;
        RECT  8.405 2.520 8.615 3.220 ;
        END
        ANTENNADIFFAREA     0.7144 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.325 0.695 11.375 1.990 ;
        RECT  11.245 0.595 11.325 1.990 ;
        RECT  11.085 0.595 11.245 3.130 ;
        RECT  11.065 0.595 11.085 1.195 ;
        RECT  10.985 2.530 11.085 3.130 ;
        END
        ANTENNADIFFAREA     0.7144 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.540 0.395 2.080 ;
        END
        ANTENNAGATEAREA     0.2236 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.700 2.470 1.990 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.835 -0.250 11.960 0.250 ;
        RECT  11.575 -0.250 11.835 1.135 ;
        RECT  10.765 -0.250 11.575 0.250 ;
        RECT  10.605 -0.250 10.765 1.135 ;
        RECT  9.730 -0.250 10.605 0.250 ;
        RECT  9.470 -0.250 9.730 0.405 ;
        RECT  8.650 -0.250 9.470 0.250 ;
        RECT  8.390 -0.250 8.650 1.220 ;
        RECT  7.570 -0.250 8.390 0.250 ;
        RECT  7.310 -0.250 7.570 0.405 ;
        RECT  4.615 -0.250 7.310 0.250 ;
        RECT  4.355 -0.250 4.615 0.405 ;
        RECT  2.095 -0.250 4.355 0.250 ;
        RECT  1.835 -0.250 2.095 0.405 ;
        RECT  0.385 -0.250 1.835 0.250 ;
        RECT  0.125 -0.250 0.385 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.755 3.440 11.960 3.940 ;
        RECT  11.495 2.265 11.755 3.940 ;
        RECT  10.735 3.440 11.495 3.940 ;
        RECT  10.475 2.605 10.735 3.940 ;
        RECT  9.330 3.440 10.475 3.940 ;
        RECT  9.070 3.285 9.330 3.940 ;
        RECT  8.195 3.440 9.070 3.940 ;
        RECT  7.935 2.605 8.195 3.940 ;
        RECT  6.655 3.440 7.935 3.940 ;
        RECT  6.395 3.285 6.655 3.940 ;
        RECT  4.035 3.440 6.395 3.940 ;
        RECT  3.775 3.285 4.035 3.940 ;
        RECT  3.015 3.440 3.775 3.940 ;
        RECT  2.755 3.285 3.015 3.940 ;
        RECT  1.955 3.440 2.755 3.940 ;
        RECT  1.695 2.990 1.955 3.940 ;
        RECT  0.385 3.440 1.695 3.940 ;
        RECT  0.125 2.475 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.385 1.735 10.545 1.995 ;
        RECT  10.060 1.735 10.385 1.900 ;
        RECT  9.900 0.935 10.060 1.900 ;
        RECT  9.835 2.505 9.935 2.765 ;
        RECT  9.835 1.740 9.900 1.900 ;
        RECT  9.675 1.740 9.835 2.765 ;
        RECT  7.965 2.180 9.675 2.340 ;
        RECT  8.855 1.380 9.115 1.980 ;
        RECT  8.155 1.420 8.855 1.580 ;
        RECT  7.995 1.075 8.155 1.580 ;
        RECT  7.850 0.635 8.110 0.895 ;
        RECT  6.905 1.075 7.995 1.235 ;
        RECT  7.705 2.180 7.965 2.380 ;
        RECT  7.030 0.655 7.850 0.815 ;
        RECT  7.025 2.335 7.185 2.920 ;
        RECT  6.770 0.470 7.030 0.815 ;
        RECT  6.905 2.335 7.025 2.495 ;
        RECT  6.675 2.760 7.025 2.920 ;
        RECT  6.745 1.075 6.905 2.495 ;
        RECT  5.120 0.470 6.770 0.630 ;
        RECT  6.150 1.075 6.745 1.235 ;
        RECT  6.515 2.760 6.675 3.080 ;
        RECT  6.395 1.680 6.555 2.580 ;
        RECT  5.490 2.920 6.515 3.080 ;
        RECT  5.800 1.680 6.395 1.840 ;
        RECT  6.335 2.420 6.395 2.580 ;
        RECT  6.175 2.420 6.335 2.735 ;
        RECT  4.415 2.575 6.175 2.735 ;
        RECT  5.985 0.820 6.150 1.235 ;
        RECT  5.880 0.820 5.985 1.080 ;
        RECT  5.825 2.130 5.985 2.395 ;
        RECT  4.925 2.130 5.825 2.290 ;
        RECT  5.540 1.385 5.800 1.840 ;
        RECT  5.370 0.820 5.630 1.085 ;
        RECT  5.165 1.680 5.540 1.840 ;
        RECT  5.225 2.920 5.490 3.130 ;
        RECT  4.585 0.925 5.370 1.085 ;
        RECT  5.005 1.265 5.165 1.840 ;
        RECT  4.960 0.470 5.120 0.745 ;
        RECT  4.860 1.265 5.005 1.425 ;
        RECT  3.595 0.585 4.960 0.745 ;
        RECT  4.825 2.130 4.925 2.395 ;
        RECT  4.665 1.750 4.825 2.395 ;
        RECT  4.585 1.750 4.665 1.910 ;
        RECT  4.425 0.925 4.585 1.910 ;
        RECT  4.105 1.295 4.425 1.455 ;
        RECT  4.300 2.125 4.415 2.735 ;
        RECT  4.140 2.125 4.300 3.105 ;
        RECT  3.985 1.655 4.245 1.915 ;
        RECT  2.395 2.945 4.140 3.105 ;
        RECT  3.845 0.965 4.105 1.455 ;
        RECT  3.805 1.755 3.985 1.915 ;
        RECT  3.465 1.295 3.845 1.455 ;
        RECT  3.645 1.755 3.805 2.765 ;
        RECT  2.555 2.605 3.645 2.765 ;
        RECT  3.335 0.495 3.595 1.095 ;
        RECT  3.305 1.295 3.465 2.425 ;
        RECT  3.075 1.295 3.305 1.455 ;
        RECT  3.205 2.165 3.305 2.425 ;
        RECT  3.010 1.690 3.110 1.850 ;
        RECT  2.975 0.655 3.075 1.455 ;
        RECT  2.850 1.690 3.010 2.330 ;
        RECT  2.815 0.655 2.975 1.500 ;
        RECT  1.155 2.170 2.850 2.330 ;
        RECT  1.625 1.340 2.815 1.500 ;
        RECT  2.465 0.880 2.565 1.140 ;
        RECT  2.295 2.510 2.555 2.765 ;
        RECT  2.305 0.585 2.465 1.140 ;
        RECT  2.135 2.945 2.395 3.260 ;
        RECT  1.545 0.585 2.305 0.745 ;
        RECT  1.515 2.605 2.295 2.765 ;
        RECT  1.385 0.430 1.545 0.745 ;
        RECT  1.355 2.605 1.515 3.055 ;
        RECT  0.735 0.430 1.385 0.590 ;
        RECT  1.205 2.815 1.355 3.055 ;
        RECT  1.105 0.915 1.205 1.175 ;
        RECT  0.735 2.815 1.205 2.975 ;
        RECT  1.105 2.035 1.155 2.635 ;
        RECT  0.945 0.915 1.105 2.635 ;
        RECT  0.575 0.430 0.735 2.975 ;
    END
END DFFSX4

MACRO DFFSX2
    CLASS CORE ;
    FOREIGN DFFSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.720 1.430 6.990 1.690 ;
        RECT  6.315 1.430 6.720 1.590 ;
        RECT  6.450 2.300 6.610 3.260 ;
        RECT  6.315 2.300 6.450 2.460 ;
        RECT  5.930 3.100 6.450 3.260 ;
        RECT  6.155 1.430 6.315 2.460 ;
        RECT  6.105 1.700 6.155 2.175 ;
        END
        ANTENNAGATEAREA     0.1456 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.835 1.390 8.995 2.340 ;
        RECT  8.635 1.390 8.835 1.550 ;
        RECT  8.575 2.180 8.835 2.340 ;
        RECT  8.475 0.470 8.635 1.550 ;
        RECT  8.415 2.180 8.575 3.220 ;
        RECT  7.830 0.470 8.475 0.630 ;
        RECT  7.720 3.060 8.415 3.220 ;
        RECT  7.570 0.470 7.830 1.110 ;
        RECT  7.560 2.390 7.720 3.220 ;
        RECT  7.460 2.390 7.560 2.995 ;
        END
        ANTENNADIFFAREA     0.6936 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.325 0.685 9.535 2.980 ;
        RECT  9.275 0.685 9.325 1.285 ;
        RECT  9.275 2.040 9.325 2.980 ;
        END
        ANTENNADIFFAREA     0.6936 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.175 0.395 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 1.490 2.335 1.650 ;
        RECT  2.075 1.490 2.235 1.990 ;
        RECT  1.965 1.700 2.075 1.990 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.975 -0.250 9.660 0.250 ;
        RECT  8.815 -0.250 8.975 1.210 ;
        RECT  7.320 -0.250 8.815 0.250 ;
        RECT  7.060 -0.250 7.320 0.855 ;
        RECT  4.105 -0.250 7.060 0.250 ;
        RECT  3.845 -0.250 4.105 0.405 ;
        RECT  2.065 -0.250 3.845 0.250 ;
        RECT  1.805 -0.250 2.065 0.405 ;
        RECT  0.385 -0.250 1.805 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.015 3.440 9.660 3.940 ;
        RECT  8.755 2.525 9.015 3.940 ;
        RECT  7.210 3.440 8.755 3.940 ;
        RECT  6.950 2.360 7.210 3.940 ;
        RECT  5.750 3.440 6.950 3.940 ;
        RECT  5.490 2.985 5.750 3.940 ;
        RECT  3.745 3.440 5.490 3.940 ;
        RECT  3.485 2.645 3.745 3.940 ;
        RECT  1.915 3.440 3.485 3.940 ;
        RECT  1.655 3.110 1.915 3.940 ;
        RECT  0.385 3.440 1.655 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.295 1.735 8.650 1.995 ;
        RECT  8.235 0.810 8.295 1.995 ;
        RECT  8.135 0.810 8.235 2.875 ;
        RECT  8.075 1.735 8.135 2.875 ;
        RECT  6.690 1.960 8.075 2.120 ;
        RECT  7.975 2.615 8.075 2.875 ;
        RECT  7.390 1.375 7.490 1.635 ;
        RECT  7.230 1.090 7.390 1.635 ;
        RECT  5.930 1.090 7.230 1.250 ;
        RECT  6.710 0.630 6.810 0.890 ;
        RECT  6.550 0.470 6.710 0.890 ;
        RECT  4.445 0.470 6.550 0.630 ;
        RECT  6.110 2.645 6.270 2.915 ;
        RECT  5.925 2.645 6.110 2.805 ;
        RECT  5.925 0.810 5.930 1.250 ;
        RECT  5.765 0.810 5.925 2.805 ;
        RECT  5.670 0.810 5.765 1.070 ;
        RECT  5.680 2.575 5.765 2.805 ;
        RECT  5.130 2.575 5.680 2.735 ;
        RECT  5.500 1.280 5.560 1.575 ;
        RECT  5.340 1.280 5.500 2.385 ;
        RECT  5.100 0.810 5.360 1.085 ;
        RECT  5.300 1.280 5.340 1.575 ;
        RECT  4.790 1.280 5.300 1.440 ;
        RECT  4.970 2.255 5.130 2.855 ;
        RECT  4.030 0.925 5.100 1.085 ;
        RECT  4.630 1.280 4.790 3.220 ;
        RECT  4.590 1.280 4.630 1.440 ;
        RECT  4.185 3.060 4.630 3.220 ;
        RECT  4.285 0.470 4.445 0.745 ;
        RECT  4.285 1.695 4.445 2.850 ;
        RECT  3.595 0.585 4.285 0.745 ;
        RECT  4.030 1.695 4.285 1.855 ;
        RECT  4.085 3.060 4.185 3.260 ;
        RECT  3.985 2.180 4.085 3.260 ;
        RECT  3.870 0.925 4.030 1.855 ;
        RECT  3.925 2.130 3.985 3.260 ;
        RECT  3.725 2.130 3.925 2.390 ;
        RECT  3.085 1.345 3.870 1.505 ;
        RECT  3.525 1.685 3.685 1.950 ;
        RECT  3.335 0.565 3.595 1.165 ;
        RECT  3.305 1.790 3.525 1.950 ;
        RECT  3.145 1.790 3.305 3.020 ;
        RECT  2.495 2.860 3.145 3.020 ;
        RECT  2.965 0.695 3.085 1.505 ;
        RECT  2.825 0.695 2.965 2.655 ;
        RECT  2.805 1.140 2.825 2.655 ;
        RECT  1.855 1.140 2.805 1.300 ;
        RECT  2.495 0.700 2.575 0.960 ;
        RECT  2.415 1.920 2.575 2.335 ;
        RECT  2.315 0.585 2.495 0.960 ;
        RECT  2.335 2.515 2.495 3.020 ;
        RECT  1.175 2.175 2.415 2.335 ;
        RECT  2.235 2.515 2.335 2.930 ;
        RECT  1.515 0.585 2.315 0.745 ;
        RECT  1.375 2.770 2.235 2.930 ;
        RECT  1.595 1.130 1.855 1.390 ;
        RECT  1.355 0.540 1.515 0.745 ;
        RECT  1.115 2.720 1.375 2.980 ;
        RECT  0.925 0.540 1.355 0.700 ;
        RECT  0.965 0.880 1.175 2.500 ;
        RECT  0.735 2.720 1.115 2.880 ;
        RECT  0.915 0.880 0.965 1.140 ;
        RECT  0.915 2.240 0.965 2.500 ;
        RECT  0.735 0.500 0.925 0.700 ;
        RECT  0.575 0.500 0.735 2.880 ;
    END
END DFFSX2

MACRO DFFSX1
    CLASS CORE ;
    FOREIGN DFFSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 1.470 6.435 1.730 ;
        RECT  6.105 1.290 6.315 1.730 ;
        RECT  6.040 1.570 6.105 1.730 ;
        RECT  5.880 1.570 6.040 3.255 ;
        RECT  5.260 3.095 5.880 3.255 ;
        END
        ANTENNAGATEAREA     0.1144 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.575 0.760 7.735 2.755 ;
        RECT  7.485 0.760 7.575 0.945 ;
        RECT  7.485 2.335 7.575 2.755 ;
        RECT  7.235 0.760 7.485 0.920 ;
        RECT  7.235 2.595 7.485 2.755 ;
        RECT  7.175 0.695 7.235 0.920 ;
        RECT  7.025 2.595 7.235 3.220 ;
        RECT  7.015 0.475 7.175 0.920 ;
        RECT  6.940 2.595 7.025 3.195 ;
        RECT  6.915 0.475 7.015 0.735 ;
        END
        ANTENNADIFFAREA     0.3796 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.090 1.105 8.155 2.585 ;
        RECT  8.075 1.105 8.090 2.750 ;
        RECT  7.915 0.920 8.075 2.750 ;
        END
        ANTENNADIFFAREA     0.3646 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.530 0.520 1.990 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 1.700 2.635 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.715 -0.250 8.280 0.250 ;
        RECT  7.455 -0.250 7.715 0.405 ;
        RECT  6.665 -0.250 7.455 0.250 ;
        RECT  6.405 -0.250 6.665 0.770 ;
        RECT  3.160 -0.250 6.405 0.250 ;
        RECT  3.000 -0.250 3.160 0.670 ;
        RECT  2.005 -0.250 3.000 0.250 ;
        RECT  1.745 -0.250 2.005 0.405 ;
        RECT  0.385 -0.250 1.745 0.250 ;
        RECT  0.125 -0.250 0.385 1.290 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.740 3.440 8.280 3.940 ;
        RECT  7.480 3.285 7.740 3.940 ;
        RECT  6.650 3.440 7.480 3.940 ;
        RECT  6.390 2.810 6.650 3.940 ;
        RECT  5.080 3.440 6.390 3.940 ;
        RECT  4.820 2.920 5.080 3.940 ;
        RECT  3.705 3.440 4.820 3.940 ;
        RECT  3.445 2.870 3.705 3.940 ;
        RECT  1.580 3.440 3.445 3.940 ;
        RECT  1.320 3.060 1.580 3.940 ;
        RECT  0.385 3.440 1.320 3.940 ;
        RECT  0.125 2.175 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.255 1.635 7.395 1.895 ;
        RECT  7.230 1.100 7.255 2.245 ;
        RECT  7.095 1.100 7.230 2.295 ;
        RECT  6.995 1.100 7.095 1.365 ;
        RECT  6.970 2.085 7.095 2.295 ;
        RECT  6.380 2.085 6.970 2.245 ;
        RECT  6.780 1.560 6.915 1.820 ;
        RECT  6.620 0.950 6.780 1.820 ;
        RECT  5.700 0.950 6.620 1.110 ;
        RECT  6.220 1.950 6.380 2.245 ;
        RECT  5.855 0.460 6.115 0.630 ;
        RECT  3.500 0.470 5.855 0.630 ;
        RECT  5.540 0.950 5.700 2.845 ;
        RECT  5.360 0.950 5.540 1.110 ;
        RECT  5.410 2.575 5.540 2.845 ;
        RECT  4.985 2.575 5.410 2.735 ;
        RECT  5.100 0.840 5.360 1.110 ;
        RECT  5.200 1.290 5.360 2.395 ;
        RECT  4.640 1.290 5.200 1.450 ;
        RECT  4.825 2.085 4.985 2.735 ;
        RECT  4.530 0.810 4.790 1.100 ;
        RECT  4.480 1.290 4.640 2.635 ;
        RECT  3.840 0.810 4.530 0.970 ;
        RECT  4.280 1.290 4.480 1.450 ;
        RECT  4.050 2.475 4.480 2.635 ;
        RECT  4.140 1.695 4.300 2.285 ;
        RECT  4.070 1.150 4.280 1.450 ;
        RECT  3.840 1.695 4.140 1.855 ;
        RECT  4.020 1.150 4.070 1.310 ;
        RECT  3.890 2.475 4.050 3.210 ;
        RECT  3.780 2.475 3.890 2.635 ;
        RECT  3.680 0.810 3.840 1.855 ;
        RECT  3.615 2.085 3.780 2.635 ;
        RECT  2.975 1.360 3.680 1.520 ;
        RECT  3.515 2.085 3.615 2.245 ;
        RECT  3.340 0.470 3.500 1.080 ;
        RECT  3.315 1.715 3.500 1.875 ;
        RECT  3.180 0.920 3.340 1.080 ;
        RECT  3.265 1.715 3.315 2.680 ;
        RECT  3.155 1.715 3.265 3.110 ;
        RECT  2.920 0.920 3.180 1.180 ;
        RECT  3.105 2.520 3.155 3.110 ;
        RECT  2.585 2.950 3.105 3.110 ;
        RECT  2.815 1.360 2.975 2.330 ;
        RECT  2.765 2.510 2.925 2.770 ;
        RECT  2.630 1.360 2.815 1.520 ;
        RECT  2.455 2.170 2.815 2.330 ;
        RECT  2.260 2.510 2.765 2.670 ;
        RECT  2.380 0.460 2.645 0.745 ;
        RECT  2.370 1.020 2.630 1.520 ;
        RECT  2.325 2.860 2.585 3.110 ;
        RECT  0.860 0.585 2.380 0.745 ;
        RECT  1.900 1.360 2.370 1.520 ;
        RECT  1.920 2.950 2.325 3.110 ;
        RECT  2.100 2.220 2.260 2.670 ;
        RECT  1.215 2.220 2.100 2.380 ;
        RECT  1.760 2.560 1.920 3.110 ;
        RECT  1.740 1.360 1.900 1.660 ;
        RECT  1.465 2.560 1.760 2.720 ;
        RECT  1.205 2.560 1.465 2.820 ;
        RECT  1.055 1.030 1.215 2.380 ;
        RECT  0.860 2.560 1.205 2.720 ;
        RECT  0.700 0.585 0.860 2.720 ;
    END
END DFFSX1

MACRO DFFSXL
    CLASS CORE ;
    FOREIGN DFFSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 1.470 6.435 1.730 ;
        RECT  6.105 1.290 6.315 1.730 ;
        RECT  6.040 1.570 6.105 1.730 ;
        RECT  5.880 1.570 6.040 3.255 ;
        RECT  5.260 3.095 5.880 3.255 ;
        END
        ANTENNAGATEAREA     0.0806 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.575 0.760 7.735 2.710 ;
        RECT  7.485 0.760 7.575 0.945 ;
        RECT  7.485 2.335 7.575 2.710 ;
        RECT  7.235 0.760 7.485 0.920 ;
        RECT  7.235 2.550 7.485 2.710 ;
        RECT  7.205 0.695 7.235 0.920 ;
        RECT  7.075 2.550 7.235 3.220 ;
        RECT  7.015 0.595 7.205 0.920 ;
        RECT  7.025 2.765 7.075 3.220 ;
        RECT  6.940 2.765 7.025 3.025 ;
        RECT  6.945 0.595 7.015 0.855 ;
        END
        ANTENNADIFFAREA     0.2238 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.095 1.105 8.155 2.175 ;
        RECT  8.090 0.920 8.095 2.175 ;
        RECT  7.930 0.920 8.090 2.575 ;
        END
        ANTENNADIFFAREA     0.2142 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.530 0.520 1.990 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 1.700 2.635 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.715 -0.250 8.280 0.250 ;
        RECT  7.455 -0.250 7.715 0.405 ;
        RECT  6.625 -0.250 7.455 0.250 ;
        RECT  6.365 -0.250 6.625 0.405 ;
        RECT  3.160 -0.250 6.365 0.250 ;
        RECT  3.000 -0.250 3.160 0.670 ;
        RECT  2.005 -0.250 3.000 0.250 ;
        RECT  1.745 -0.250 2.005 0.405 ;
        RECT  0.385 -0.250 1.745 0.250 ;
        RECT  0.125 -0.250 0.385 1.290 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.740 3.440 8.280 3.940 ;
        RECT  7.480 2.895 7.740 3.940 ;
        RECT  6.650 3.440 7.480 3.940 ;
        RECT  6.390 2.810 6.650 3.940 ;
        RECT  5.080 3.440 6.390 3.940 ;
        RECT  4.820 3.035 5.080 3.940 ;
        RECT  3.705 3.440 4.820 3.940 ;
        RECT  3.445 3.035 3.705 3.940 ;
        RECT  1.580 3.440 3.445 3.940 ;
        RECT  1.320 3.115 1.580 3.940 ;
        RECT  0.385 3.440 1.320 3.940 ;
        RECT  0.125 2.175 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.255 1.635 7.395 1.895 ;
        RECT  7.095 1.100 7.255 2.345 ;
        RECT  6.995 1.100 7.095 1.365 ;
        RECT  6.970 2.085 7.095 2.345 ;
        RECT  6.380 2.085 6.970 2.245 ;
        RECT  6.780 1.560 6.915 1.820 ;
        RECT  6.620 0.950 6.780 1.820 ;
        RECT  5.700 0.950 6.620 1.110 ;
        RECT  6.220 1.950 6.380 2.245 ;
        RECT  5.855 0.460 6.115 0.630 ;
        RECT  3.500 0.470 5.855 0.630 ;
        RECT  5.540 0.950 5.700 2.845 ;
        RECT  5.360 0.950 5.540 1.110 ;
        RECT  4.985 2.685 5.540 2.845 ;
        RECT  5.100 0.840 5.360 1.110 ;
        RECT  5.200 1.290 5.360 2.395 ;
        RECT  4.640 1.290 5.200 1.450 ;
        RECT  4.825 2.025 4.985 2.845 ;
        RECT  4.530 0.810 4.790 1.100 ;
        RECT  4.480 1.290 4.640 2.635 ;
        RECT  3.840 0.810 4.530 0.970 ;
        RECT  4.280 1.290 4.480 1.450 ;
        RECT  4.045 2.475 4.480 2.635 ;
        RECT  4.130 1.695 4.290 2.285 ;
        RECT  4.070 1.150 4.280 1.450 ;
        RECT  3.840 1.695 4.130 1.855 ;
        RECT  4.020 1.150 4.070 1.310 ;
        RECT  3.885 2.475 4.045 3.260 ;
        RECT  3.780 2.475 3.885 2.635 ;
        RECT  3.680 0.810 3.840 1.855 ;
        RECT  3.615 2.085 3.780 2.635 ;
        RECT  2.975 1.360 3.680 1.520 ;
        RECT  3.515 2.085 3.615 2.245 ;
        RECT  3.340 0.470 3.500 1.080 ;
        RECT  3.315 1.700 3.500 1.860 ;
        RECT  3.215 0.920 3.340 1.080 ;
        RECT  3.265 1.700 3.315 2.680 ;
        RECT  3.155 1.700 3.265 3.110 ;
        RECT  2.955 0.920 3.215 1.180 ;
        RECT  3.105 2.520 3.155 3.110 ;
        RECT  2.585 2.950 3.105 3.110 ;
        RECT  2.815 1.360 2.975 2.330 ;
        RECT  2.765 2.510 2.925 2.770 ;
        RECT  2.630 1.360 2.815 1.520 ;
        RECT  2.455 2.170 2.815 2.330 ;
        RECT  2.260 2.510 2.765 2.670 ;
        RECT  2.380 0.460 2.645 0.745 ;
        RECT  2.370 0.930 2.630 1.520 ;
        RECT  2.325 2.860 2.585 3.110 ;
        RECT  0.860 0.585 2.380 0.745 ;
        RECT  1.900 1.360 2.370 1.520 ;
        RECT  1.920 2.950 2.325 3.110 ;
        RECT  2.100 2.220 2.260 2.670 ;
        RECT  1.215 2.220 2.100 2.380 ;
        RECT  1.760 2.560 1.920 3.110 ;
        RECT  1.740 1.360 1.900 1.660 ;
        RECT  1.465 2.560 1.760 2.720 ;
        RECT  1.205 2.560 1.465 2.820 ;
        RECT  1.055 1.030 1.215 2.380 ;
        RECT  0.860 2.560 1.205 2.720 ;
        RECT  0.700 0.585 0.860 2.720 ;
    END
END DFFSXL

MACRO DFFRX4
    CLASS CORE ;
    FOREIGN DFFRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.890 1.460 9.530 1.620 ;
        RECT  8.820 1.290 8.890 1.620 ;
        RECT  8.660 0.470 8.820 1.620 ;
        RECT  5.670 0.470 8.660 0.630 ;
        RECT  5.660 0.470 5.670 0.760 ;
        RECT  5.500 0.470 5.660 1.040 ;
        RECT  5.395 0.880 5.500 1.040 ;
        RECT  5.370 0.880 5.395 1.170 ;
        RECT  5.030 0.880 5.370 1.380 ;
        RECT  4.960 0.880 5.030 1.040 ;
        RECT  4.800 0.470 4.960 1.040 ;
        RECT  3.375 0.470 4.800 0.630 ;
        RECT  3.215 0.470 3.375 0.745 ;
        RECT  2.105 0.585 3.215 0.745 ;
        RECT  1.945 0.585 2.105 1.380 ;
        RECT  1.770 1.220 1.945 1.380 ;
        RECT  1.610 1.220 1.770 1.605 ;
        RECT  1.510 1.345 1.610 1.605 ;
        END
        ANTENNAGATEAREA     0.3510 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.115 0.620 11.135 1.220 ;
        RECT  10.960 0.620 11.115 1.555 ;
        RECT  10.875 0.620 10.960 2.755 ;
        RECT  10.720 1.105 10.875 2.755 ;
        RECT  10.705 1.105 10.720 2.175 ;
        END
        ANTENNADIFFAREA     0.8312 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.155 1.090 12.330 2.400 ;
        RECT  12.090 0.675 12.155 2.400 ;
        RECT  11.895 0.675 12.090 1.330 ;
        RECT  12.085 1.515 12.090 2.400 ;
        RECT  12.080 2.045 12.085 2.400 ;
        RECT  11.820 2.155 12.080 3.095 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.175 1.550 0.440 2.030 ;
        RECT  0.125 1.700 0.175 1.990 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.575 2.470 1.925 ;
        RECT  2.135 1.575 2.175 1.990 ;
        RECT  1.965 1.700 2.135 1.990 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.665 -0.250 12.880 0.250 ;
        RECT  12.405 -0.250 12.665 0.865 ;
        RECT  11.645 -0.250 12.405 0.250 ;
        RECT  11.385 -0.250 11.645 1.170 ;
        RECT  10.590 -0.250 11.385 0.250 ;
        RECT  10.330 -0.250 10.590 0.405 ;
        RECT  9.280 -0.250 10.330 0.250 ;
        RECT  9.020 -0.250 9.280 0.405 ;
        RECT  5.300 -0.250 9.020 0.250 ;
        RECT  5.140 -0.250 5.300 0.625 ;
        RECT  2.990 -0.250 5.140 0.250 ;
        RECT  2.050 -0.250 2.990 0.405 ;
        RECT  0.000 -0.250 2.050 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.630 3.440 12.880 3.940 ;
        RECT  12.370 2.605 12.630 3.940 ;
        RECT  11.510 3.405 12.370 3.940 ;
        RECT  11.250 3.285 11.510 3.940 ;
        RECT  10.400 3.405 11.250 3.940 ;
        RECT  10.140 3.285 10.400 3.940 ;
        RECT  9.230 3.405 10.140 3.940 ;
        RECT  8.970 3.285 9.230 3.940 ;
        RECT  6.445 3.405 8.970 3.940 ;
        RECT  6.185 2.975 6.445 3.940 ;
        RECT  5.110 3.440 6.185 3.940 ;
        RECT  4.950 2.560 5.110 3.940 ;
        RECT  4.575 3.440 4.950 3.940 ;
        RECT  4.315 2.800 4.575 3.940 ;
        RECT  2.760 3.440 4.315 3.940 ;
        RECT  2.500 3.285 2.760 3.940 ;
        RECT  0.395 3.440 2.500 3.940 ;
        RECT  0.135 2.275 0.395 3.940 ;
        RECT  0.000 3.440 0.135 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.645 1.585 11.905 1.845 ;
        RECT  11.435 1.685 11.645 1.845 ;
        RECT  11.275 1.685 11.435 3.100 ;
        RECT  10.395 2.940 11.275 3.100 ;
        RECT  10.235 0.915 10.395 3.100 ;
        RECT  10.180 0.915 10.235 1.975 ;
        RECT  9.820 2.910 10.235 3.100 ;
        RECT  10.165 0.695 10.180 1.975 ;
        RECT  9.920 0.695 10.165 1.295 ;
        RECT  8.690 1.815 10.165 1.975 ;
        RECT  9.795 2.155 10.055 2.415 ;
        RECT  9.560 2.595 9.820 3.195 ;
        RECT  8.480 2.155 9.795 2.315 ;
        RECT  6.890 3.020 8.655 3.180 ;
        RECT  8.320 0.810 8.480 2.825 ;
        RECT  7.480 0.810 8.320 0.970 ;
        RECT  8.185 2.155 8.320 2.825 ;
        RECT  7.430 2.600 8.185 2.825 ;
        RECT  7.890 1.150 8.020 1.310 ;
        RECT  7.890 2.255 7.940 2.415 ;
        RECT  7.730 1.150 7.890 2.415 ;
        RECT  6.010 1.700 7.730 1.860 ;
        RECT  7.680 2.255 7.730 2.415 ;
        RECT  7.270 0.810 7.480 1.230 ;
        RECT  7.170 2.205 7.430 2.825 ;
        RECT  7.220 0.970 7.270 1.230 ;
        RECT  6.870 0.880 6.970 1.140 ;
        RECT  5.845 2.285 6.920 2.445 ;
        RECT  6.730 2.625 6.890 3.180 ;
        RECT  6.710 0.880 6.870 1.345 ;
        RECT  5.455 2.625 6.730 2.785 ;
        RECT  6.010 1.185 6.710 1.345 ;
        RECT  5.850 1.135 6.010 1.860 ;
        RECT  5.845 1.700 5.850 1.860 ;
        RECT  5.685 1.700 5.845 2.445 ;
        RECT  4.965 1.700 5.685 1.865 ;
        RECT  5.635 2.285 5.685 2.445 ;
        RECT  5.295 2.090 5.455 2.785 ;
        RECT  4.620 2.090 5.295 2.250 ;
        RECT  4.805 1.650 4.965 1.910 ;
        RECT  4.225 2.430 4.735 2.590 ;
        RECT  4.460 0.810 4.620 2.250 ;
        RECT  3.770 0.810 4.460 0.970 ;
        RECT  4.225 1.150 4.275 1.310 ;
        RECT  4.065 1.150 4.225 2.590 ;
        RECT  4.015 1.150 4.065 1.310 ;
        RECT  3.685 2.425 4.065 2.590 ;
        RECT  3.770 1.555 3.830 1.815 ;
        RECT  3.730 0.810 3.770 1.815 ;
        RECT  3.610 0.810 3.730 2.160 ;
        RECT  3.525 2.425 3.685 3.080 ;
        RECT  3.385 0.970 3.610 1.230 ;
        RECT  3.570 1.555 3.610 2.160 ;
        RECT  3.260 2.000 3.570 2.160 ;
        RECT  3.475 2.430 3.525 3.080 ;
        RECT  3.425 2.720 3.475 3.080 ;
        RECT  1.330 2.920 3.425 3.080 ;
        RECT  3.065 1.450 3.320 1.710 ;
        RECT  3.240 2.000 3.260 2.295 ;
        RECT  3.080 2.000 3.240 2.735 ;
        RECT  1.445 2.575 3.080 2.735 ;
        RECT  2.905 1.030 3.065 1.710 ;
        RECT  2.545 1.030 2.905 1.190 ;
        RECT  2.835 1.550 2.905 1.710 ;
        RECT  2.675 1.550 2.835 2.385 ;
        RECT  1.785 2.225 2.675 2.385 ;
        RECT  2.285 0.930 2.545 1.190 ;
        RECT  1.625 1.790 1.785 2.385 ;
        RECT  1.375 0.475 1.635 0.735 ;
        RECT  1.235 1.790 1.625 1.950 ;
        RECT  1.285 2.130 1.445 2.735 ;
        RECT  0.385 0.575 1.375 0.735 ;
        RECT  1.070 2.920 1.330 3.200 ;
        RECT  1.235 1.415 1.285 1.575 ;
        RECT  1.075 1.415 1.235 1.950 ;
        RECT  0.950 0.975 1.210 1.235 ;
        RECT  1.025 1.415 1.075 1.575 ;
        RECT  0.800 2.920 1.070 3.080 ;
        RECT  0.800 1.075 0.950 1.235 ;
        RECT  0.640 1.075 0.800 3.080 ;
        RECT  0.125 0.560 0.385 1.160 ;
    END
END DFFRX4

MACRO DFFRX2
    CLASS CORE ;
    FOREIGN DFFRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.160 1.435 7.255 1.695 ;
        RECT  6.995 1.430 7.160 1.695 ;
        RECT  6.610 1.430 6.995 1.590 ;
        RECT  6.450 0.470 6.610 1.590 ;
        RECT  5.335 0.470 6.450 0.630 ;
        RECT  5.175 0.470 5.335 1.380 ;
        RECT  4.655 1.220 5.175 1.380 ;
        RECT  4.495 0.470 4.655 1.380 ;
        RECT  3.170 0.470 4.495 0.630 ;
        RECT  3.010 0.470 3.170 0.745 ;
        RECT  1.715 0.585 3.010 0.745 ;
        RECT  1.555 0.585 1.715 1.170 ;
        RECT  1.535 0.880 1.555 1.170 ;
        RECT  1.505 0.880 1.535 1.660 ;
        RECT  1.375 0.945 1.505 1.660 ;
        END
        ANTENNAGATEAREA     0.2080 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.590 1.515 8.615 2.175 ;
        RECT  8.470 1.515 8.590 2.755 ;
        RECT  8.330 0.515 8.470 2.755 ;
        RECT  8.310 0.515 8.330 1.925 ;
        RECT  8.180 0.515 8.310 0.775 ;
        END
        ANTENNADIFFAREA     0.4844 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.350 2.155 9.565 2.755 ;
        RECT  9.360 0.845 9.460 1.105 ;
        RECT  9.200 0.845 9.360 1.450 ;
        RECT  9.305 2.110 9.350 2.755 ;
        RECT  9.165 2.110 9.305 2.315 ;
        RECT  9.165 1.290 9.200 1.450 ;
        RECT  9.005 1.290 9.165 2.315 ;
        RECT  8.865 1.290 9.005 1.765 ;
        END
        ANTENNADIFFAREA     0.4028 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.585 0.845 1.845 ;
        RECT  0.765 1.585 0.795 1.990 ;
        RECT  0.495 1.585 0.765 2.040 ;
        END
        ANTENNAGATEAREA     0.1313 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 1.310 2.280 1.570 ;
        RECT  2.175 1.310 2.230 1.650 ;
        RECT  1.965 1.290 2.175 1.650 ;
        RECT  1.775 1.420 1.965 1.650 ;
        END
        ANTENNAGATEAREA     0.0650 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.970 -0.250 10.120 0.250 ;
        RECT  9.710 -0.250 9.970 1.095 ;
        RECT  9.010 -0.250 9.710 0.250 ;
        RECT  8.750 -0.250 9.010 1.040 ;
        RECT  7.155 -0.250 8.750 0.250 ;
        RECT  8.690 0.780 8.750 1.040 ;
        RECT  6.895 -0.250 7.155 1.140 ;
        RECT  4.995 -0.250 6.895 0.250 ;
        RECT  4.835 -0.250 4.995 0.625 ;
        RECT  2.805 -0.250 4.835 0.250 ;
        RECT  2.545 -0.250 2.805 0.405 ;
        RECT  1.705 -0.250 2.545 0.250 ;
        RECT  1.445 -0.250 1.705 0.405 ;
        RECT  0.000 -0.250 1.445 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.965 3.440 10.120 3.940 ;
        RECT  9.705 3.285 9.965 3.940 ;
        RECT  8.990 3.440 9.705 3.940 ;
        RECT  8.390 3.285 8.990 3.940 ;
        RECT  6.875 3.440 8.390 3.940 ;
        RECT  6.615 3.285 6.875 3.940 ;
        RECT  4.805 3.440 6.615 3.940 ;
        RECT  4.645 2.560 4.805 3.940 ;
        RECT  4.270 3.440 4.645 3.940 ;
        RECT  4.010 2.800 4.270 3.940 ;
        RECT  2.510 3.440 4.010 3.940 ;
        RECT  2.250 3.285 2.510 3.940 ;
        RECT  0.555 3.440 2.250 3.940 ;
        RECT  0.295 3.285 0.555 3.940 ;
        RECT  0.000 3.440 0.295 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.800 1.725 9.960 3.105 ;
        RECT  9.735 1.725 9.800 1.885 ;
        RECT  8.075 2.945 9.800 3.105 ;
        RECT  9.475 1.625 9.735 1.885 ;
        RECT  8.025 1.885 8.075 3.105 ;
        RECT  8.020 1.035 8.025 3.105 ;
        RECT  7.860 1.035 8.020 3.110 ;
        RECT  7.765 1.035 7.860 2.045 ;
        RECT  7.445 2.950 7.860 3.110 ;
        RECT  6.755 1.885 7.765 2.045 ;
        RECT  7.420 2.305 7.680 2.565 ;
        RECT  7.185 2.950 7.445 3.210 ;
        RECT  6.215 2.400 7.420 2.560 ;
        RECT  6.495 1.785 6.755 2.045 ;
        RECT  6.020 2.980 6.280 3.240 ;
        RECT  6.215 0.820 6.265 0.980 ;
        RECT  6.075 0.820 6.215 2.560 ;
        RECT  6.055 0.820 6.075 2.780 ;
        RECT  6.005 0.820 6.055 0.980 ;
        RECT  5.815 2.180 6.055 2.780 ;
        RECT  5.160 3.030 6.020 3.190 ;
        RECT  5.545 0.820 5.705 1.860 ;
        RECT  5.515 1.700 5.545 1.860 ;
        RECT  5.355 1.700 5.515 2.770 ;
        RECT  4.660 1.700 5.355 1.860 ;
        RECT  5.000 2.090 5.160 3.190 ;
        RECT  4.315 2.090 5.000 2.250 ;
        RECT  4.500 1.650 4.660 1.910 ;
        RECT  3.870 2.430 4.430 2.590 ;
        RECT  4.155 0.810 4.315 2.250 ;
        RECT  3.525 0.810 4.155 0.970 ;
        RECT  3.870 1.150 3.970 1.310 ;
        RECT  3.710 1.150 3.870 2.590 ;
        RECT  3.330 2.430 3.710 2.590 ;
        RECT  3.365 0.810 3.525 1.105 ;
        RECT  3.230 1.555 3.450 1.815 ;
        RECT  3.330 0.945 3.365 1.105 ;
        RECT  3.230 0.945 3.330 1.205 ;
        RECT  3.170 2.430 3.330 3.050 ;
        RECT  3.070 0.945 3.230 2.230 ;
        RECT  0.310 2.890 3.170 3.050 ;
        RECT  2.985 2.070 3.070 2.230 ;
        RECT  2.825 2.070 2.985 2.645 ;
        RECT  1.245 2.485 2.825 2.645 ;
        RECT  2.640 1.630 2.820 1.890 ;
        RECT  2.480 0.950 2.640 2.180 ;
        RECT  1.965 0.950 2.480 1.110 ;
        RECT  2.080 2.020 2.480 2.180 ;
        RECT  1.980 2.020 2.080 2.280 ;
        RECT  1.820 1.840 1.980 2.280 ;
        RECT  1.185 1.840 1.820 2.000 ;
        RECT  1.085 2.200 1.245 2.645 ;
        RECT  1.025 1.140 1.185 2.000 ;
        RECT  0.985 2.200 1.085 2.360 ;
        RECT  0.650 1.140 1.025 1.300 ;
        RECT  0.490 1.040 0.650 1.300 ;
        RECT  0.310 0.570 0.530 0.830 ;
        RECT  0.270 0.570 0.310 3.050 ;
        RECT  0.150 0.620 0.270 3.050 ;
    END
END DFFRX2

MACRO DFFRX1
    CLASS CORE ;
    FOREIGN DFFRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.430 6.845 1.795 ;
        RECT  6.585 1.290 6.775 1.795 ;
        RECT  6.565 1.290 6.585 1.600 ;
        RECT  6.315 1.430 6.565 1.600 ;
        RECT  6.205 1.105 6.315 1.600 ;
        RECT  6.035 0.470 6.205 1.600 ;
        RECT  4.885 0.470 6.035 0.640 ;
        RECT  4.715 0.470 4.885 1.335 ;
        RECT  4.525 1.165 4.715 1.335 ;
        RECT  4.265 1.165 4.525 1.430 ;
        RECT  4.195 1.165 4.265 1.325 ;
        RECT  4.035 0.470 4.195 1.325 ;
        RECT  2.725 0.470 4.035 0.630 ;
        RECT  2.565 0.470 2.725 0.745 ;
        RECT  1.530 0.585 2.565 0.745 ;
        RECT  1.420 0.585 1.530 0.760 ;
        RECT  1.260 0.585 1.420 1.075 ;
        END
        ANTENNAGATEAREA     0.1274 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.960 1.700 8.155 1.990 ;
        RECT  7.800 0.690 7.960 2.315 ;
        RECT  7.590 0.690 7.800 0.850 ;
        RECT  7.670 2.110 7.800 2.315 ;
        RECT  7.640 2.155 7.670 2.315 ;
        RECT  7.380 2.155 7.640 2.755 ;
        RECT  7.330 0.565 7.590 0.850 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 0.845 8.615 2.755 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.640 0.885 1.900 ;
        RECT  0.585 1.640 0.835 2.100 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.385 1.995 1.645 ;
        RECT  1.505 1.290 1.715 1.645 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.160 -0.250 8.740 0.250 ;
        RECT  7.900 -0.250 8.160 0.405 ;
        RECT  6.670 -0.250 7.900 0.250 ;
        RECT  6.410 -0.250 6.670 0.405 ;
        RECT  4.535 -0.250 6.410 0.250 ;
        RECT  4.375 -0.250 4.535 0.625 ;
        RECT  2.365 -0.250 4.375 0.250 ;
        RECT  2.105 -0.250 2.365 0.405 ;
        RECT  0.000 -0.250 2.105 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.040 3.440 8.740 3.940 ;
        RECT  7.440 3.285 8.040 3.940 ;
        RECT  6.055 3.440 7.440 3.940 ;
        RECT  5.795 3.285 6.055 3.940 ;
        RECT  3.810 3.440 5.795 3.940 ;
        RECT  3.550 2.800 3.810 3.940 ;
        RECT  2.320 3.440 3.550 3.940 ;
        RECT  1.720 3.285 2.320 3.940 ;
        RECT  0.410 3.440 1.720 3.940 ;
        RECT  0.150 3.285 0.410 3.940 ;
        RECT  0.000 3.440 0.150 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.200 2.945 8.445 3.105 ;
        RECT  7.285 1.130 7.545 1.390 ;
        RECT  7.200 1.180 7.285 1.390 ;
        RECT  7.040 1.180 7.200 3.130 ;
        RECT  6.210 1.980 7.040 2.140 ;
        RECT  6.625 2.970 7.040 3.130 ;
        RECT  6.600 2.550 6.860 2.790 ;
        RECT  6.365 2.970 6.625 3.230 ;
        RECT  5.750 2.550 6.600 2.710 ;
        RECT  5.950 1.785 6.210 2.140 ;
        RECT  5.750 0.820 5.850 0.980 ;
        RECT  5.590 0.820 5.750 2.710 ;
        RECT  5.285 2.500 5.590 2.710 ;
        RECT  4.275 3.030 5.485 3.190 ;
        RECT  5.025 2.500 5.285 2.760 ;
        RECT  5.070 0.830 5.230 1.860 ;
        RECT  4.615 1.700 5.070 1.860 ;
        RECT  4.615 2.495 4.715 2.755 ;
        RECT  4.455 1.700 4.615 2.755 ;
        RECT  4.200 1.700 4.455 1.860 ;
        RECT  4.115 2.090 4.275 3.190 ;
        RECT  4.040 1.650 4.200 1.910 ;
        RECT  3.855 2.090 4.115 2.250 ;
        RECT  3.515 2.430 3.905 2.590 ;
        RECT  3.695 0.810 3.855 2.250 ;
        RECT  3.070 0.810 3.695 0.970 ;
        RECT  3.355 1.150 3.515 2.590 ;
        RECT  3.250 1.150 3.355 1.310 ;
        RECT  3.310 2.430 3.355 2.590 ;
        RECT  3.150 2.430 3.310 2.950 ;
        RECT  0.290 2.790 3.150 2.950 ;
        RECT  3.070 1.540 3.115 1.800 ;
        RECT  3.015 0.810 3.070 1.800 ;
        RECT  2.910 0.810 3.015 2.185 ;
        RECT  2.735 0.980 2.910 1.240 ;
        RECT  2.865 1.540 2.910 2.185 ;
        RECT  2.855 1.540 2.865 2.575 ;
        RECT  2.705 2.025 2.855 2.575 ;
        RECT  0.950 2.415 2.705 2.575 ;
        RECT  2.525 1.585 2.595 1.845 ;
        RECT  2.495 0.950 2.525 1.845 ;
        RECT  2.365 0.950 2.495 2.100 ;
        RECT  1.670 0.950 2.365 1.110 ;
        RECT  2.335 1.585 2.365 2.100 ;
        RECT  1.795 1.940 2.335 2.100 ;
        RECT  1.535 1.940 1.795 2.230 ;
        RECT  1.275 1.940 1.535 2.100 ;
        RECT  1.115 1.260 1.275 2.100 ;
        RECT  0.630 1.260 1.115 1.420 ;
        RECT  0.690 2.355 0.950 2.575 ;
        RECT  0.470 1.020 0.630 1.420 ;
        RECT  0.290 0.490 0.480 0.750 ;
        RECT  0.220 0.490 0.290 2.950 ;
        RECT  0.130 0.540 0.220 2.950 ;
    END
END DFFRX1

MACRO DFFRXL
    CLASS CORE ;
    FOREIGN DFFRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.475 6.845 1.745 ;
        RECT  6.585 1.290 6.775 1.745 ;
        RECT  6.565 1.290 6.585 1.645 ;
        RECT  6.315 1.475 6.565 1.645 ;
        RECT  6.205 1.105 6.315 1.645 ;
        RECT  6.035 0.470 6.205 1.645 ;
        RECT  4.885 0.470 6.035 0.640 ;
        RECT  4.715 0.470 4.885 1.335 ;
        RECT  4.525 1.165 4.715 1.335 ;
        RECT  4.265 1.165 4.525 1.430 ;
        RECT  4.195 1.165 4.265 1.325 ;
        RECT  4.035 0.470 4.195 1.325 ;
        RECT  2.690 0.470 4.035 0.630 ;
        RECT  2.530 0.470 2.690 0.745 ;
        RECT  1.420 0.585 2.530 0.745 ;
        RECT  1.260 0.585 1.420 1.075 ;
        END
        ANTENNAGATEAREA     0.1001 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.960 1.700 8.155 1.990 ;
        RECT  7.800 0.690 7.960 2.315 ;
        RECT  7.560 0.690 7.800 0.850 ;
        RECT  7.670 2.110 7.800 2.315 ;
        RECT  7.640 2.155 7.670 2.315 ;
        RECT  7.480 2.155 7.640 2.585 ;
        RECT  7.300 0.565 7.560 0.850 ;
        RECT  7.380 2.325 7.480 2.585 ;
        END
        ANTENNADIFFAREA     0.2135 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 0.845 8.615 2.585 ;
        END
        ANTENNADIFFAREA     0.2135 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.690 0.885 1.950 ;
        RECT  0.585 1.690 0.835 2.150 ;
        END
        ANTENNAGATEAREA     0.0442 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.385 1.995 1.645 ;
        RECT  1.505 1.290 1.715 1.645 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.160 -0.250 8.740 0.250 ;
        RECT  7.900 -0.250 8.160 0.405 ;
        RECT  6.670 -0.250 7.900 0.250 ;
        RECT  6.410 -0.250 6.670 0.405 ;
        RECT  4.535 -0.250 6.410 0.250 ;
        RECT  4.375 -0.250 4.535 0.625 ;
        RECT  2.340 -0.250 4.375 0.250 ;
        RECT  2.080 -0.250 2.340 0.405 ;
        RECT  1.680 -0.250 2.080 0.250 ;
        RECT  1.420 -0.250 1.680 0.405 ;
        RECT  0.000 -0.250 1.420 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.040 3.440 8.740 3.940 ;
        RECT  7.440 3.285 8.040 3.940 ;
        RECT  6.055 3.440 7.440 3.940 ;
        RECT  5.795 3.285 6.055 3.940 ;
        RECT  3.810 3.440 5.795 3.940 ;
        RECT  3.550 2.800 3.810 3.940 ;
        RECT  2.325 3.440 3.550 3.940 ;
        RECT  1.725 3.285 2.325 3.940 ;
        RECT  0.410 3.440 1.725 3.940 ;
        RECT  0.150 3.285 0.410 3.940 ;
        RECT  0.000 3.440 0.150 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.220 2.895 8.480 3.155 ;
        RECT  7.200 2.895 8.220 3.055 ;
        RECT  7.285 1.130 7.545 1.390 ;
        RECT  7.200 1.180 7.285 1.390 ;
        RECT  7.040 1.180 7.200 3.160 ;
        RECT  6.210 1.935 7.040 2.095 ;
        RECT  6.365 3.000 7.040 3.160 ;
        RECT  6.600 2.550 6.860 2.790 ;
        RECT  5.750 2.550 6.600 2.710 ;
        RECT  5.950 1.835 6.210 2.095 ;
        RECT  5.750 0.820 5.850 0.980 ;
        RECT  5.590 0.820 5.750 2.710 ;
        RECT  5.285 2.500 5.590 2.710 ;
        RECT  4.245 3.030 5.485 3.190 ;
        RECT  5.025 2.500 5.285 2.760 ;
        RECT  5.070 0.830 5.230 1.860 ;
        RECT  4.615 1.700 5.070 1.860 ;
        RECT  4.615 2.495 4.715 2.755 ;
        RECT  4.455 1.700 4.615 2.755 ;
        RECT  4.200 1.700 4.455 1.860 ;
        RECT  4.085 2.090 4.245 3.190 ;
        RECT  4.040 1.650 4.200 1.910 ;
        RECT  3.855 2.090 4.085 2.250 ;
        RECT  3.515 2.430 3.905 2.590 ;
        RECT  3.695 0.810 3.855 2.250 ;
        RECT  3.070 0.810 3.695 0.970 ;
        RECT  3.355 1.150 3.515 2.590 ;
        RECT  3.250 1.150 3.355 1.310 ;
        RECT  3.310 2.430 3.355 2.590 ;
        RECT  3.150 2.430 3.310 2.950 ;
        RECT  0.285 2.790 3.150 2.950 ;
        RECT  3.070 1.540 3.115 1.800 ;
        RECT  3.015 0.810 3.070 1.800 ;
        RECT  2.910 0.810 3.015 2.185 ;
        RECT  2.705 0.945 2.910 1.205 ;
        RECT  2.865 1.540 2.910 2.185 ;
        RECT  2.855 1.540 2.865 2.575 ;
        RECT  2.705 2.025 2.855 2.575 ;
        RECT  0.690 2.415 2.705 2.575 ;
        RECT  2.495 1.450 2.595 1.710 ;
        RECT  2.335 0.945 2.495 2.100 ;
        RECT  1.640 0.945 2.335 1.105 ;
        RECT  1.795 1.940 2.335 2.100 ;
        RECT  1.535 1.940 1.795 2.230 ;
        RECT  1.275 1.940 1.535 2.100 ;
        RECT  1.115 1.260 1.275 2.100 ;
        RECT  0.630 1.260 1.115 1.420 ;
        RECT  0.470 1.020 0.630 1.420 ;
        RECT  0.285 0.525 0.480 0.785 ;
        RECT  0.220 0.525 0.285 2.950 ;
        RECT  0.125 0.575 0.220 2.950 ;
    END
END DFFRXL

MACRO DFFQXL
    CLASS CORE ;
    FOREIGN DFFQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 0.585 6.785 2.710 ;
        RECT  6.625 0.585 6.775 2.810 ;
        RECT  6.545 0.585 6.625 0.945 ;
        RECT  6.565 1.760 6.625 2.810 ;
        RECT  6.130 2.550 6.565 2.810 ;
        END
        ANTENNADIFFAREA     0.2569 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.530 0.395 1.995 ;
        END
        ANTENNAGATEAREA     0.0507 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.955 1.700 3.095 1.990 ;
        RECT  2.695 1.700 2.955 2.135 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.810 -0.250 6.900 0.250 ;
        RECT  5.210 -0.250 5.810 0.595 ;
        RECT  3.670 -0.250 5.210 0.250 ;
        RECT  3.410 -0.250 3.670 0.405 ;
        RECT  2.095 -0.250 3.410 0.250 ;
        RECT  1.935 -0.250 2.095 0.675 ;
        RECT  0.385 -0.250 1.935 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.415 3.440 6.900 3.940 ;
        RECT  5.475 3.285 6.415 3.940 ;
        RECT  4.190 3.440 5.475 3.940 ;
        RECT  3.930 3.285 4.190 3.940 ;
        RECT  2.285 3.440 3.930 3.940 ;
        RECT  1.685 3.055 2.285 3.940 ;
        RECT  0.385 3.440 1.685 3.940 ;
        RECT  0.125 2.500 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.345 1.225 6.445 1.485 ;
        RECT  6.185 0.775 6.345 1.485 ;
        RECT  5.765 2.025 6.230 2.285 ;
        RECT  5.300 0.775 6.185 0.935 ;
        RECT  5.765 1.155 6.005 1.315 ;
        RECT  5.605 1.155 5.765 2.955 ;
        RECT  5.245 2.795 5.605 2.955 ;
        RECT  5.140 0.775 5.300 2.615 ;
        RECT  5.085 2.795 5.245 3.230 ;
        RECT  4.305 0.775 5.140 0.960 ;
        RECT  4.735 2.455 5.140 2.615 ;
        RECT  4.795 1.140 4.955 2.270 ;
        RECT  4.060 0.430 4.825 0.590 ;
        RECT  4.060 1.140 4.795 1.300 ;
        RECT  4.395 2.110 4.795 2.270 ;
        RECT  4.575 2.455 4.735 2.800 ;
        RECT  4.325 1.575 4.585 1.840 ;
        RECT  4.235 2.110 4.395 3.105 ;
        RECT  3.435 1.575 4.325 1.735 ;
        RECT  2.995 2.945 4.235 3.105 ;
        RECT  3.900 0.430 4.060 1.300 ;
        RECT  3.895 1.915 4.055 2.765 ;
        RECT  3.435 0.585 3.900 0.745 ;
        RECT  3.025 2.605 3.895 2.765 ;
        RECT  3.175 0.585 3.435 0.775 ;
        RECT  3.275 1.160 3.435 2.425 ;
        RECT  3.235 1.160 3.275 1.320 ;
        RECT  3.210 2.165 3.275 2.425 ;
        RECT  2.975 0.955 3.235 1.320 ;
        RECT  2.715 0.585 3.175 0.745 ;
        RECT  2.865 2.375 3.025 2.765 ;
        RECT  2.735 2.945 2.995 3.205 ;
        RECT  1.755 0.955 2.975 1.115 ;
        RECT  2.515 2.375 2.865 2.535 ;
        RECT  2.685 2.945 2.735 3.105 ;
        RECT  2.455 0.465 2.715 0.745 ;
        RECT  2.525 2.715 2.685 3.105 ;
        RECT  2.515 1.295 2.650 1.455 ;
        RECT  1.240 2.715 2.525 2.875 ;
        RECT  2.355 1.295 2.515 2.535 ;
        RECT  1.675 2.375 2.355 2.535 ;
        RECT  2.015 1.545 2.175 1.875 ;
        RECT  1.415 1.715 2.015 1.875 ;
        RECT  1.595 0.535 1.755 1.115 ;
        RECT  1.515 2.105 1.675 2.535 ;
        RECT  1.435 0.535 1.595 0.695 ;
        RECT  1.415 2.105 1.515 2.265 ;
        RECT  1.175 0.435 1.435 0.695 ;
        RECT  1.255 0.875 1.415 1.875 ;
        RECT  0.735 0.875 1.255 1.035 ;
        RECT  1.235 2.715 1.240 3.125 ;
        RECT  1.075 2.055 1.235 3.125 ;
        RECT  0.915 1.265 1.075 2.215 ;
        RECT  0.935 2.865 1.075 3.125 ;
        RECT  0.735 2.525 0.895 2.685 ;
        RECT  0.575 0.875 0.735 2.685 ;
    END
END DFFQXL

MACRO DFFQX4
    CLASS CORE ;
    FOREIGN DFFQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.405 0.620 8.530 1.220 ;
        RECT  8.270 0.620 8.405 3.140 ;
        RECT  8.145 0.880 8.270 3.140 ;
        RECT  7.945 0.880 8.145 1.580 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.115 1.330 0.395 1.995 ;
        END
        ANTENNAGATEAREA     0.1092 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.530 3.095 1.990 ;
        RECT  2.750 1.700 2.885 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.040 -0.250 9.200 0.250 ;
        RECT  8.780 -0.250 9.040 1.100 ;
        RECT  7.905 -0.250 8.780 0.250 ;
        RECT  6.965 -0.250 7.905 0.615 ;
        RECT  5.505 -0.250 6.965 0.250 ;
        RECT  5.245 -0.250 5.505 0.405 ;
        RECT  4.145 -0.250 5.245 0.250 ;
        RECT  3.885 -0.250 4.145 0.405 ;
        RECT  2.805 -0.250 3.885 0.250 ;
        RECT  2.545 -0.250 2.805 0.405 ;
        RECT  0.385 -0.250 2.545 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.945 3.440 9.200 3.940 ;
        RECT  8.685 2.200 8.945 3.940 ;
        RECT  7.735 3.440 8.685 3.940 ;
        RECT  7.475 2.895 7.735 3.940 ;
        RECT  6.795 3.005 7.475 3.940 ;
        RECT  5.410 3.440 6.795 3.940 ;
        RECT  5.150 3.285 5.410 3.940 ;
        RECT  4.050 3.440 5.150 3.940 ;
        RECT  3.790 3.285 4.050 3.940 ;
        RECT  2.815 3.440 3.790 3.940 ;
        RECT  2.555 3.285 2.815 3.940 ;
        RECT  1.885 3.440 2.555 3.940 ;
        RECT  1.625 3.285 1.885 3.940 ;
        RECT  0.385 3.440 1.625 3.940 ;
        RECT  0.125 2.775 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.465 1.035 7.625 2.270 ;
        RECT  7.410 1.035 7.465 1.295 ;
        RECT  7.125 2.010 7.465 2.270 ;
        RECT  6.785 1.475 7.285 1.735 ;
        RECT  6.965 2.010 7.125 2.780 ;
        RECT  6.410 2.620 6.965 2.780 ;
        RECT  6.625 0.575 6.785 2.440 ;
        RECT  6.385 0.575 6.625 0.735 ;
        RECT  6.210 2.280 6.625 2.440 ;
        RECT  6.210 3.100 6.520 3.260 ;
        RECT  6.385 1.255 6.445 1.515 ;
        RECT  6.125 0.455 6.385 0.745 ;
        RECT  6.225 0.925 6.385 2.100 ;
        RECT  4.085 0.925 6.225 1.085 ;
        RECT  5.870 1.940 6.225 2.100 ;
        RECT  6.050 2.280 6.210 2.710 ;
        RECT  6.050 2.945 6.210 3.260 ;
        RECT  4.395 0.585 6.125 0.745 ;
        RECT  4.560 2.285 6.050 2.445 ;
        RECT  4.115 2.945 6.050 3.105 ;
        RECT  5.910 1.580 6.010 1.740 ;
        RECT  5.750 1.265 5.910 1.740 ;
        RECT  5.710 1.940 5.870 2.105 ;
        RECT  3.745 1.265 5.750 1.425 ;
        RECT  4.115 1.945 5.710 2.105 ;
        RECT  3.775 1.605 5.350 1.765 ;
        RECT  4.300 2.285 4.560 2.545 ;
        RECT  3.955 1.945 4.115 3.105 ;
        RECT  3.925 0.605 4.085 1.085 ;
        RECT  3.385 2.945 3.955 3.105 ;
        RECT  3.345 0.605 3.925 0.765 ;
        RECT  3.615 1.605 3.775 2.685 ;
        RECT  3.485 1.005 3.745 1.425 ;
        RECT  2.515 2.525 3.615 2.685 ;
        RECT  3.435 1.155 3.485 1.425 ;
        RECT  3.275 1.155 3.435 2.185 ;
        RECT  3.125 2.945 3.385 3.215 ;
        RECT  3.085 0.495 3.345 0.765 ;
        RECT  2.895 1.155 3.275 1.315 ;
        RECT  1.365 2.945 3.125 3.105 ;
        RECT  2.735 0.905 2.895 1.315 ;
        RECT  1.755 0.905 2.735 1.065 ;
        RECT  2.515 1.245 2.545 1.505 ;
        RECT  2.355 1.245 2.515 2.685 ;
        RECT  2.285 1.245 2.355 1.505 ;
        RECT  2.185 2.325 2.355 2.585 ;
        RECT  1.675 2.325 2.185 2.485 ;
        RECT  2.015 1.715 2.175 1.975 ;
        RECT  1.415 1.715 2.015 1.875 ;
        RECT  1.595 0.580 1.755 1.065 ;
        RECT  1.515 2.100 1.675 2.485 ;
        RECT  1.435 0.580 1.595 0.740 ;
        RECT  1.415 2.100 1.515 2.260 ;
        RECT  1.175 0.475 1.435 0.740 ;
        RECT  1.255 0.920 1.415 1.875 ;
        RECT  1.235 2.945 1.365 3.260 ;
        RECT  0.735 0.920 1.255 1.080 ;
        RECT  1.105 2.055 1.235 3.260 ;
        RECT  1.075 2.055 1.105 3.105 ;
        RECT  0.915 1.260 1.075 2.215 ;
        RECT  0.735 2.735 0.895 2.995 ;
        RECT  0.575 0.920 0.735 2.895 ;
    END
END DFFQX4

MACRO DFFQX2
    CLASS CORE ;
    FOREIGN DFFQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.195 2.200 7.235 2.995 ;
        RECT  7.050 2.200 7.195 3.140 ;
        RECT  6.955 2.110 7.050 3.140 ;
        RECT  6.935 0.620 6.955 3.140 ;
        RECT  6.765 0.620 6.935 2.700 ;
        RECT  6.600 0.620 6.765 1.220 ;
        RECT  6.590 0.620 6.600 1.170 ;
        RECT  6.565 0.690 6.590 1.170 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.530 0.395 1.995 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.530 3.095 1.990 ;
        RECT  2.695 1.700 2.885 1.990 ;
        END
        ANTENNAGATEAREA     0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.150 -0.250 7.360 0.250 ;
        RECT  5.210 -0.250 6.150 0.565 ;
        RECT  3.670 -0.250 5.210 0.250 ;
        RECT  3.410 -0.250 3.670 0.405 ;
        RECT  2.340 -0.250 3.410 0.250 ;
        RECT  2.080 -0.250 2.340 0.775 ;
        RECT  0.385 -0.250 2.080 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.355 3.440 7.360 3.940 ;
        RECT  5.415 2.945 6.355 3.940 ;
        RECT  3.865 3.440 5.415 3.940 ;
        RECT  3.605 3.285 3.865 3.940 ;
        RECT  1.885 3.440 3.605 3.940 ;
        RECT  1.625 3.285 1.885 3.940 ;
        RECT  0.385 3.440 1.625 3.940 ;
        RECT  0.125 2.520 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.285 1.475 6.385 1.735 ;
        RECT  6.125 0.745 6.285 1.735 ;
        RECT  5.915 2.010 6.265 2.270 ;
        RECT  5.300 0.745 6.125 0.905 ;
        RECT  5.830 1.085 5.945 1.245 ;
        RECT  5.830 2.010 5.915 2.765 ;
        RECT  5.670 1.085 5.830 2.765 ;
        RECT  5.005 2.605 5.670 2.765 ;
        RECT  5.140 0.745 5.300 2.315 ;
        RECT  4.295 0.770 5.140 0.930 ;
        RECT  4.715 2.155 5.140 2.315 ;
        RECT  4.720 2.945 4.980 3.260 ;
        RECT  4.795 1.110 4.955 1.975 ;
        RECT  4.115 0.430 4.935 0.590 ;
        RECT  4.115 1.110 4.795 1.270 ;
        RECT  4.265 1.815 4.795 1.975 ;
        RECT  4.265 2.945 4.720 3.105 ;
        RECT  4.455 2.155 4.715 2.755 ;
        RECT  4.145 1.460 4.405 1.635 ;
        RECT  4.105 1.815 4.265 3.105 ;
        RECT  3.435 1.460 4.145 1.620 ;
        RECT  3.955 0.430 4.115 1.270 ;
        RECT  3.355 2.945 4.105 3.105 ;
        RECT  3.435 0.585 3.955 0.745 ;
        RECT  3.780 1.800 3.925 1.960 ;
        RECT  3.620 1.800 3.780 2.720 ;
        RECT  2.835 2.560 3.620 2.720 ;
        RECT  3.175 0.585 3.435 0.785 ;
        RECT  3.275 1.190 3.435 2.375 ;
        RECT  3.095 2.945 3.355 3.215 ;
        RECT  3.220 1.190 3.275 1.350 ;
        RECT  3.015 2.215 3.275 2.375 ;
        RECT  2.995 1.090 3.220 1.350 ;
        RECT  2.925 0.585 3.175 0.775 ;
        RECT  2.495 2.945 3.095 3.105 ;
        RECT  2.835 0.955 2.995 1.350 ;
        RECT  2.665 0.515 2.925 0.775 ;
        RECT  1.755 0.955 2.835 1.115 ;
        RECT  2.675 2.375 2.835 2.720 ;
        RECT  2.515 2.375 2.675 2.535 ;
        RECT  2.515 1.295 2.650 1.455 ;
        RECT  2.355 1.295 2.515 2.535 ;
        RECT  2.335 2.715 2.495 3.105 ;
        RECT  1.675 2.375 2.355 2.535 ;
        RECT  1.235 2.715 2.335 2.875 ;
        RECT  2.015 1.715 2.175 1.975 ;
        RECT  1.415 1.715 2.015 1.875 ;
        RECT  1.595 0.535 1.755 1.115 ;
        RECT  1.515 2.105 1.675 2.535 ;
        RECT  1.435 0.535 1.595 0.695 ;
        RECT  1.415 2.105 1.515 2.265 ;
        RECT  1.175 0.435 1.435 0.695 ;
        RECT  1.255 0.925 1.415 1.875 ;
        RECT  0.735 0.925 1.255 1.085 ;
        RECT  1.075 2.055 1.235 3.165 ;
        RECT  0.915 1.265 1.075 2.215 ;
        RECT  0.935 2.905 1.075 3.165 ;
        RECT  0.735 2.565 0.895 2.725 ;
        RECT  0.575 0.925 0.735 2.725 ;
    END
END DFFQX2

MACRO DFFQX1
    CLASS CORE ;
    FOREIGN DFFQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 0.475 6.785 2.700 ;
        RECT  6.625 0.475 6.775 2.810 ;
        RECT  6.545 0.475 6.625 0.735 ;
        RECT  6.565 1.925 6.625 2.810 ;
        RECT  6.315 2.540 6.565 2.810 ;
        RECT  6.310 2.540 6.315 2.800 ;
        END
        ANTENNADIFFAREA     0.3764 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.530 0.395 1.995 ;
        END
        ANTENNAGATEAREA     0.0507 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.955 1.700 3.095 1.990 ;
        RECT  2.695 1.700 2.955 2.135 ;
        END
        ANTENNAGATEAREA     0.0806 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.810 -0.250 6.900 0.250 ;
        RECT  5.210 -0.250 5.810 0.595 ;
        RECT  3.670 -0.250 5.210 0.250 ;
        RECT  3.410 -0.250 3.670 0.405 ;
        RECT  2.095 -0.250 3.410 0.250 ;
        RECT  1.935 -0.250 2.095 0.735 ;
        RECT  0.385 -0.250 1.935 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.415 3.440 6.900 3.940 ;
        RECT  5.475 3.285 6.415 3.940 ;
        RECT  3.850 3.440 5.475 3.940 ;
        RECT  3.590 3.285 3.850 3.940 ;
        RECT  2.285 3.440 3.590 3.940 ;
        RECT  1.685 3.055 2.285 3.940 ;
        RECT  0.385 3.440 1.685 3.940 ;
        RECT  0.125 2.500 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.345 1.225 6.445 1.485 ;
        RECT  6.185 0.775 6.345 1.485 ;
        RECT  5.765 2.025 6.230 2.285 ;
        RECT  5.300 0.775 6.185 0.935 ;
        RECT  5.765 1.155 6.005 1.315 ;
        RECT  5.605 1.155 5.765 2.955 ;
        RECT  5.245 2.795 5.605 2.955 ;
        RECT  5.140 0.775 5.300 2.615 ;
        RECT  5.085 2.795 5.245 3.230 ;
        RECT  4.305 0.775 5.140 0.960 ;
        RECT  4.735 2.455 5.140 2.615 ;
        RECT  4.795 1.140 4.955 2.270 ;
        RECT  4.060 0.430 4.825 0.590 ;
        RECT  4.060 1.140 4.795 1.300 ;
        RECT  4.395 2.110 4.795 2.270 ;
        RECT  4.575 2.455 4.735 3.065 ;
        RECT  4.325 1.570 4.585 1.830 ;
        RECT  4.235 2.110 4.395 3.105 ;
        RECT  3.435 1.570 4.325 1.730 ;
        RECT  2.965 2.945 4.235 3.105 ;
        RECT  3.900 0.430 4.060 1.300 ;
        RECT  3.895 1.915 4.055 2.175 ;
        RECT  3.435 0.585 3.900 0.745 ;
        RECT  3.800 2.015 3.895 2.175 ;
        RECT  3.640 2.015 3.800 2.765 ;
        RECT  3.025 2.605 3.640 2.765 ;
        RECT  3.175 0.585 3.435 0.775 ;
        RECT  3.275 1.160 3.435 2.425 ;
        RECT  3.235 1.160 3.275 1.320 ;
        RECT  3.210 2.165 3.275 2.425 ;
        RECT  2.975 0.955 3.235 1.320 ;
        RECT  2.715 0.585 3.175 0.745 ;
        RECT  2.865 2.375 3.025 2.765 ;
        RECT  1.755 0.955 2.975 1.115 ;
        RECT  2.705 2.945 2.965 3.215 ;
        RECT  2.515 2.375 2.865 2.535 ;
        RECT  2.455 0.465 2.715 0.745 ;
        RECT  2.685 2.945 2.705 3.105 ;
        RECT  2.525 2.715 2.685 3.105 ;
        RECT  2.515 1.295 2.650 1.455 ;
        RECT  1.240 2.715 2.525 2.875 ;
        RECT  2.355 1.295 2.515 2.535 ;
        RECT  1.675 2.375 2.355 2.535 ;
        RECT  2.015 1.545 2.175 1.875 ;
        RECT  1.415 1.715 2.015 1.875 ;
        RECT  1.595 0.535 1.755 1.115 ;
        RECT  1.515 2.105 1.675 2.535 ;
        RECT  1.435 0.535 1.595 0.695 ;
        RECT  1.415 2.105 1.515 2.265 ;
        RECT  1.175 0.435 1.435 0.695 ;
        RECT  1.255 0.875 1.415 1.875 ;
        RECT  0.735 0.875 1.255 1.035 ;
        RECT  1.235 2.715 1.240 3.125 ;
        RECT  1.075 2.055 1.235 3.125 ;
        RECT  0.915 1.265 1.075 2.215 ;
        RECT  0.935 2.865 1.075 3.125 ;
        RECT  0.735 2.525 0.895 2.685 ;
        RECT  0.575 0.875 0.735 2.685 ;
    END
END DFFQX1

MACRO DFFX4
    CLASS CORE ;
    FOREIGN DFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.845 1.035 10.915 2.585 ;
        RECT  10.655 0.695 10.845 2.895 ;
        RECT  10.585 0.695 10.655 1.295 ;
        RECT  10.585 1.955 10.655 2.895 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.825 1.515 9.995 1.765 ;
        RECT  9.565 0.695 9.825 2.215 ;
        RECT  9.325 1.290 9.565 1.990 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.850 0.795 2.400 ;
        RECT  0.535 1.850 0.585 2.175 ;
        END
        ANTENNAGATEAREA     0.1274 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.685 1.895 2.945 2.155 ;
        RECT  2.635 1.995 2.685 2.155 ;
        RECT  2.475 1.995 2.635 2.400 ;
        RECT  2.425 2.110 2.475 2.400 ;
        END
        ANTENNAGATEAREA     0.2002 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 -0.250 11.500 0.250 ;
        RECT  11.095 -0.250 11.355 1.095 ;
        RECT  10.335 -0.250 11.095 0.250 ;
        RECT  10.075 -0.250 10.335 1.095 ;
        RECT  9.315 -0.250 10.075 0.250 ;
        RECT  9.055 -0.250 9.315 0.755 ;
        RECT  8.400 -0.250 9.055 0.250 ;
        RECT  8.155 -0.250 8.400 1.250 ;
        RECT  8.085 -0.250 8.155 0.405 ;
        RECT  6.525 -0.250 8.085 0.250 ;
        RECT  6.265 -0.250 6.525 0.575 ;
        RECT  4.855 -0.250 6.265 0.250 ;
        RECT  4.595 -0.250 4.855 0.895 ;
        RECT  3.165 -0.250 4.595 0.250 ;
        RECT  2.905 -0.250 3.165 0.745 ;
        RECT  2.255 -0.250 2.905 0.250 ;
        RECT  1.995 -0.250 2.255 0.945 ;
        RECT  0.485 -0.250 1.995 0.250 ;
        RECT  0.225 -0.250 0.485 1.065 ;
        RECT  0.000 -0.250 0.225 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 3.440 11.500 3.940 ;
        RECT  11.095 2.255 11.355 3.940 ;
        RECT  10.335 3.440 11.095 3.940 ;
        RECT  10.075 2.935 10.335 3.940 ;
        RECT  9.315 3.440 10.075 3.940 ;
        RECT  9.055 2.935 9.315 3.940 ;
        RECT  8.375 3.440 9.055 3.940 ;
        RECT  8.115 2.545 8.375 3.940 ;
        RECT  6.525 3.440 8.115 3.940 ;
        RECT  6.265 2.715 6.525 3.940 ;
        RECT  4.825 3.440 6.265 3.940 ;
        RECT  4.565 3.285 4.825 3.940 ;
        RECT  3.325 3.440 4.565 3.940 ;
        RECT  3.065 3.285 3.325 3.940 ;
        RECT  2.265 3.440 3.065 3.940 ;
        RECT  2.005 3.285 2.265 3.940 ;
        RECT  0.625 3.440 2.005 3.940 ;
        RECT  0.365 2.580 0.625 3.940 ;
        RECT  0.000 3.440 0.365 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.375 1.515 10.475 1.775 ;
        RECT  10.215 1.515 10.375 2.585 ;
        RECT  8.915 2.425 10.215 2.585 ;
        RECT  8.865 1.035 8.915 1.295 ;
        RECT  8.865 1.985 8.915 2.585 ;
        RECT  8.705 1.035 8.865 2.585 ;
        RECT  8.655 1.035 8.705 1.295 ;
        RECT  8.655 1.980 8.705 2.585 ;
        RECT  7.885 1.980 8.655 2.140 ;
        RECT  8.265 1.515 8.525 1.775 ;
        RECT  7.975 1.565 8.265 1.775 ;
        RECT  7.815 0.755 7.975 1.775 ;
        RECT  7.885 2.855 7.935 3.115 ;
        RECT  7.725 1.980 7.885 3.115 ;
        RECT  7.375 0.755 7.815 0.915 ;
        RECT  7.545 1.615 7.815 1.775 ;
        RECT  7.675 2.855 7.725 3.115 ;
        RECT  7.205 1.145 7.635 1.405 ;
        RECT  7.385 1.615 7.545 2.535 ;
        RECT  7.375 2.375 7.385 2.535 ;
        RECT  7.115 0.705 7.375 0.965 ;
        RECT  7.115 2.375 7.375 2.990 ;
        RECT  7.045 1.145 7.205 2.195 ;
        RECT  5.415 0.755 7.115 0.915 ;
        RECT  5.675 2.375 7.115 2.535 ;
        RECT  6.670 1.145 7.045 1.305 ;
        RECT  6.945 1.805 7.045 2.195 ;
        RECT  5.365 1.805 6.945 1.965 ;
        RECT  6.510 1.095 6.670 1.305 ;
        RECT  4.685 1.095 6.510 1.255 ;
        RECT  5.025 1.435 6.325 1.595 ;
        RECT  5.415 2.375 5.675 2.975 ;
        RECT  5.205 1.805 5.365 2.170 ;
        RECT  4.915 2.010 5.205 2.170 ;
        RECT  4.865 1.435 5.025 1.830 ;
        RECT  4.755 2.010 4.915 3.105 ;
        RECT  4.535 1.670 4.865 1.830 ;
        RECT  1.135 2.945 4.755 3.105 ;
        RECT  4.525 1.095 4.685 1.390 ;
        RECT  4.375 1.670 4.535 2.765 ;
        RECT  4.515 1.230 4.525 1.390 ;
        RECT  4.255 1.230 4.515 1.490 ;
        RECT  3.675 2.605 4.375 2.765 ;
        RECT  4.075 0.790 4.345 1.050 ;
        RECT  4.075 2.045 4.125 2.305 ;
        RECT  3.915 0.470 4.075 2.305 ;
        RECT  3.725 0.470 3.915 0.630 ;
        RECT  3.865 2.045 3.915 2.305 ;
        RECT  3.675 0.825 3.725 1.085 ;
        RECT  3.515 0.825 3.675 2.765 ;
        RECT  3.465 0.825 3.515 1.085 ;
        RECT  2.205 2.605 3.515 2.765 ;
        RECT  3.220 1.265 3.320 1.525 ;
        RECT  3.060 1.265 3.220 1.715 ;
        RECT  1.475 1.555 3.060 1.715 ;
        RECT  2.505 0.995 2.765 1.285 ;
        RECT  1.815 1.125 2.505 1.285 ;
        RECT  2.045 1.915 2.205 2.765 ;
        RECT  1.945 1.915 2.045 2.175 ;
        RECT  1.655 0.545 1.815 1.285 ;
        RECT  0.930 0.545 1.655 0.705 ;
        RECT  1.315 0.895 1.475 2.625 ;
        RECT  1.115 0.895 1.315 1.155 ;
        RECT  0.975 1.355 1.135 3.105 ;
        RECT  0.930 1.355 0.975 1.620 ;
        RECT  0.770 0.545 0.930 1.620 ;
    END
END DFFX4

MACRO DFFX2
    CLASS CORE ;
    FOREIGN DFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.405 0.695 8.615 3.045 ;
        RECT  8.355 0.695 8.405 1.295 ;
        RECT  8.355 2.105 8.405 3.045 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.060 1.700 7.235 1.990 ;
        RECT  7.050 0.495 7.215 0.755 ;
        RECT  6.930 1.700 7.060 2.215 ;
        RECT  6.955 0.495 7.050 0.760 ;
        RECT  6.930 0.595 6.955 0.760 ;
        RECT  6.770 0.595 6.930 2.215 ;
        END
        ANTENNADIFFAREA     0.6173 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.530 0.460 1.990 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 2.110 2.755 2.400 ;
        END
        ANTENNAGATEAREA     0.1144 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.075 -0.250 8.740 0.250 ;
        RECT  7.815 -0.250 8.075 0.645 ;
        RECT  6.670 -0.250 7.815 0.250 ;
        RECT  6.410 -0.250 6.670 0.405 ;
        RECT  4.520 -0.250 6.410 0.250 ;
        RECT  4.260 -0.250 4.520 0.635 ;
        RECT  3.120 -0.250 4.260 0.250 ;
        RECT  2.180 -0.250 3.120 0.405 ;
        RECT  0.400 -0.250 2.180 0.250 ;
        RECT  0.140 -0.250 0.400 0.405 ;
        RECT  0.000 -0.250 0.140 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.075 3.440 8.740 3.940 ;
        RECT  7.815 2.205 8.075 3.940 ;
        RECT  6.510 3.440 7.815 3.940 ;
        RECT  6.250 2.890 6.510 3.940 ;
        RECT  4.320 3.440 6.250 3.940 ;
        RECT  4.060 3.285 4.320 3.940 ;
        RECT  3.300 3.440 4.060 3.940 ;
        RECT  3.040 3.285 3.300 3.940 ;
        RECT  2.240 3.440 3.040 3.940 ;
        RECT  1.980 3.285 2.240 3.940 ;
        RECT  0.650 3.440 1.980 3.940 ;
        RECT  0.390 2.170 0.650 3.940 ;
        RECT  0.000 3.440 0.390 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.615 1.585 8.215 1.845 ;
        RECT  7.455 1.035 7.615 2.725 ;
        RECT  7.355 1.035 7.455 1.295 ;
        RECT  7.265 2.465 7.455 2.725 ;
        RECT  6.070 2.465 7.265 2.625 ;
        RECT  6.340 0.610 6.500 2.130 ;
        RECT  6.230 0.610 6.340 0.770 ;
        RECT  5.725 1.970 6.340 2.130 ;
        RECT  6.070 0.470 6.230 0.770 ;
        RECT  5.940 0.950 6.100 1.790 ;
        RECT  5.450 0.470 6.070 0.630 ;
        RECT  5.910 2.465 6.070 2.905 ;
        RECT  5.890 0.950 5.940 1.110 ;
        RECT  5.385 1.630 5.940 1.790 ;
        RECT  5.810 2.645 5.910 2.905 ;
        RECT  5.680 0.810 5.890 1.110 ;
        RECT  5.020 1.290 5.760 1.450 ;
        RECT  5.565 1.970 5.725 2.455 ;
        RECT  5.630 0.810 5.680 1.075 ;
        RECT  4.330 0.915 5.630 1.075 ;
        RECT  5.175 2.295 5.565 2.455 ;
        RECT  5.290 0.470 5.450 0.735 ;
        RECT  5.225 1.630 5.385 2.115 ;
        RECT  4.670 1.955 5.225 2.115 ;
        RECT  4.915 2.295 5.175 2.895 ;
        RECT  4.860 1.275 5.020 1.450 ;
        RECT  3.990 1.275 4.860 1.435 ;
        RECT  4.510 1.955 4.670 3.105 ;
        RECT  2.750 2.945 4.510 3.105 ;
        RECT  4.330 1.615 4.430 1.775 ;
        RECT  4.170 0.815 4.330 1.075 ;
        RECT  4.170 1.615 4.330 2.735 ;
        RECT  3.240 2.575 4.170 2.735 ;
        RECT  3.830 0.595 3.990 2.225 ;
        RECT  3.700 0.595 3.830 0.755 ;
        RECT  3.730 2.015 3.830 2.225 ;
        RECT  3.470 2.015 3.730 2.275 ;
        RECT  3.440 0.495 3.700 0.755 ;
        RECT  3.490 1.015 3.650 1.645 ;
        RECT  3.240 1.485 3.490 1.645 ;
        RECT  1.940 0.590 3.440 0.750 ;
        RECT  3.080 1.485 3.240 2.735 ;
        RECT  1.990 1.770 3.080 1.930 ;
        RECT  1.450 1.430 2.900 1.590 ;
        RECT  1.600 1.060 2.760 1.220 ;
        RECT  2.490 2.595 2.750 3.105 ;
        RECT  1.700 2.945 2.490 3.105 ;
        RECT  1.730 1.770 1.990 2.030 ;
        RECT  1.780 0.470 1.940 0.750 ;
        RECT  1.440 2.915 1.700 3.175 ;
        RECT  1.440 0.670 1.600 1.220 ;
        RECT  1.290 1.430 1.450 2.430 ;
        RECT  0.920 0.670 1.440 0.830 ;
        RECT  1.110 2.965 1.440 3.125 ;
        RECT  1.260 1.430 1.290 1.590 ;
        RECT  1.100 1.010 1.260 1.590 ;
        RECT  0.950 1.810 1.110 3.125 ;
        RECT  0.920 1.810 0.950 1.970 ;
        RECT  0.760 0.670 0.920 1.970 ;
        RECT  0.730 1.380 0.760 1.640 ;
    END
END DFFX2

MACRO DFFX1
    CLASS CORE ;
    FOREIGN DFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.215 2.520 7.235 2.915 ;
        RECT  7.055 0.970 7.215 2.915 ;
        RECT  7.050 0.970 7.055 1.355 ;
        RECT  7.025 2.520 7.055 2.915 ;
        RECT  6.955 0.970 7.050 1.230 ;
        RECT  6.975 2.655 7.025 2.915 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.765 1.425 6.870 2.425 ;
        RECT  6.710 0.695 6.765 2.425 ;
        RECT  6.605 0.695 6.710 1.585 ;
        RECT  6.320 2.265 6.710 2.425 ;
        RECT  6.035 0.695 6.605 0.855 ;
        RECT  6.315 2.265 6.320 2.745 ;
        RECT  6.265 2.265 6.315 2.995 ;
        RECT  6.105 2.265 6.265 3.225 ;
        RECT  5.975 2.965 6.105 3.225 ;
        RECT  5.775 0.540 6.035 0.855 ;
        END
        ANTENNADIFFAREA     0.3300 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.955 0.385 2.535 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.805 1.605 3.095 2.055 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.620 -0.250 7.360 0.250 ;
        RECT  6.360 -0.250 6.620 0.405 ;
        RECT  5.470 -0.250 6.360 0.250 ;
        RECT  5.210 -0.250 5.470 0.405 ;
        RECT  3.735 -0.250 5.210 0.250 ;
        RECT  3.475 -0.250 3.735 0.405 ;
        RECT  2.105 -0.250 3.475 0.250 ;
        RECT  1.945 -0.250 2.105 0.735 ;
        RECT  0.385 -0.250 1.945 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.805 3.440 7.360 3.940 ;
        RECT  6.545 3.285 6.805 3.940 ;
        RECT  5.385 3.440 6.545 3.940 ;
        RECT  5.125 3.285 5.385 3.940 ;
        RECT  3.625 3.440 5.125 3.940 ;
        RECT  3.365 3.285 3.625 3.940 ;
        RECT  1.975 3.440 3.365 3.940 ;
        RECT  1.715 3.285 1.975 3.940 ;
        RECT  0.385 3.440 1.715 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.425 1.775 6.530 2.035 ;
        RECT  6.265 1.145 6.425 2.085 ;
        RECT  5.685 1.145 6.265 1.305 ;
        RECT  5.765 1.925 6.265 2.085 ;
        RECT  5.790 1.485 6.050 1.745 ;
        RECT  5.765 2.455 5.865 2.715 ;
        RECT  5.130 1.485 5.790 1.645 ;
        RECT  5.605 1.925 5.765 2.715 ;
        RECT  5.570 1.925 5.605 2.085 ;
        RECT  5.410 1.825 5.570 2.085 ;
        RECT  5.310 1.825 5.410 1.985 ;
        RECT  4.970 0.790 5.130 2.505 ;
        RECT  4.260 0.790 4.970 0.950 ;
        RECT  4.455 2.345 4.970 2.505 ;
        RECT  4.630 1.135 4.790 2.065 ;
        RECT  4.530 1.135 4.630 1.325 ;
        RECT  4.315 1.905 4.630 2.065 ;
        RECT  3.775 1.135 4.530 1.295 ;
        RECT  4.295 2.345 4.455 2.705 ;
        RECT  4.115 1.905 4.315 2.165 ;
        RECT  3.435 1.475 4.310 1.635 ;
        RECT  3.955 1.905 4.115 3.105 ;
        RECT  1.545 2.945 3.955 3.105 ;
        RECT  3.615 0.585 3.775 1.295 ;
        RECT  3.615 1.870 3.775 2.765 ;
        RECT  2.975 0.585 3.615 0.745 ;
        RECT  2.455 2.605 3.615 2.765 ;
        RECT  3.275 1.095 3.435 2.425 ;
        RECT  3.155 1.095 3.275 1.255 ;
        RECT  2.825 2.265 3.275 2.425 ;
        RECT  2.895 0.925 3.155 1.255 ;
        RECT  2.815 0.495 2.975 0.745 ;
        RECT  1.750 0.925 2.895 1.085 ;
        RECT  2.465 0.495 2.815 0.655 ;
        RECT  2.455 1.265 2.595 2.215 ;
        RECT  2.435 1.265 2.455 2.765 ;
        RECT  2.325 1.265 2.435 1.425 ;
        RECT  2.295 2.055 2.435 2.765 ;
        RECT  2.195 2.055 2.295 2.555 ;
        RECT  1.995 1.615 2.255 1.875 ;
        RECT  1.775 2.055 2.195 2.215 ;
        RECT  1.410 1.615 1.995 1.775 ;
        RECT  1.515 1.955 1.775 2.215 ;
        RECT  1.590 0.460 1.750 1.085 ;
        RECT  1.135 0.460 1.590 0.620 ;
        RECT  1.385 2.425 1.545 3.105 ;
        RECT  1.250 0.830 1.410 1.775 ;
        RECT  1.295 2.425 1.385 2.585 ;
        RECT  1.135 1.955 1.295 2.585 ;
        RECT  0.525 0.830 1.250 0.990 ;
        RECT  0.945 2.845 1.205 3.105 ;
        RECT  1.070 1.955 1.135 2.215 ;
        RECT  1.035 1.200 1.070 2.215 ;
        RECT  0.910 1.200 1.035 2.125 ;
        RECT  0.725 2.845 0.945 3.005 ;
        RECT  0.735 1.200 0.910 1.360 ;
        RECT  0.565 1.615 0.725 3.005 ;
        RECT  0.525 1.615 0.565 1.775 ;
        RECT  0.365 0.830 0.525 1.775 ;
    END
END DFFX1

MACRO DFFXL
    CLASS CORE ;
    FOREIGN DFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.075 0.970 7.235 2.915 ;
        RECT  7.050 0.970 7.075 1.355 ;
        RECT  7.025 2.520 7.075 2.915 ;
        RECT  6.975 0.970 7.050 1.230 ;
        RECT  6.975 2.655 7.025 2.915 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.425 6.870 2.425 ;
        RECT  6.710 1.105 6.775 2.425 ;
        RECT  6.680 1.105 6.710 1.585 ;
        RECT  6.320 2.265 6.710 2.425 ;
        RECT  6.520 0.695 6.680 1.585 ;
        RECT  6.005 0.695 6.520 0.855 ;
        RECT  6.315 2.265 6.320 2.745 ;
        RECT  6.265 2.265 6.315 2.995 ;
        RECT  6.105 2.265 6.265 3.225 ;
        RECT  5.975 2.965 6.105 3.225 ;
        RECT  5.745 0.540 6.005 0.855 ;
        END
        ANTENNADIFFAREA     0.2304 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.955 0.385 2.535 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.805 1.605 3.095 2.055 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.620 -0.250 7.360 0.250 ;
        RECT  6.360 -0.250 6.620 0.405 ;
        RECT  5.470 -0.250 6.360 0.250 ;
        RECT  5.210 -0.250 5.470 0.405 ;
        RECT  3.735 -0.250 5.210 0.250 ;
        RECT  3.475 -0.250 3.735 0.405 ;
        RECT  2.105 -0.250 3.475 0.250 ;
        RECT  1.945 -0.250 2.105 0.735 ;
        RECT  0.385 -0.250 1.945 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.805 3.440 7.360 3.940 ;
        RECT  6.545 3.285 6.805 3.940 ;
        RECT  5.385 3.440 6.545 3.940 ;
        RECT  5.125 3.285 5.385 3.940 ;
        RECT  3.625 3.440 5.125 3.940 ;
        RECT  3.365 3.285 3.625 3.940 ;
        RECT  1.975 3.440 3.365 3.940 ;
        RECT  1.715 3.285 1.975 3.940 ;
        RECT  0.385 3.440 1.715 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.340 1.775 6.530 2.085 ;
        RECT  6.180 1.145 6.340 2.085 ;
        RECT  5.685 1.145 6.180 1.305 ;
        RECT  5.815 1.925 6.180 2.085 ;
        RECT  5.840 1.485 6.000 1.745 ;
        RECT  5.130 1.485 5.840 1.645 ;
        RECT  5.655 1.925 5.815 2.715 ;
        RECT  5.570 1.925 5.655 2.085 ;
        RECT  5.410 1.825 5.570 2.085 ;
        RECT  5.310 1.825 5.410 1.985 ;
        RECT  4.970 0.790 5.130 2.505 ;
        RECT  4.260 0.790 4.970 0.950 ;
        RECT  4.455 2.345 4.970 2.505 ;
        RECT  4.630 1.135 4.790 2.065 ;
        RECT  4.530 1.135 4.630 1.325 ;
        RECT  4.315 1.905 4.630 2.065 ;
        RECT  3.775 1.135 4.530 1.295 ;
        RECT  4.295 2.345 4.455 2.605 ;
        RECT  4.115 1.905 4.315 2.165 ;
        RECT  3.435 1.475 4.310 1.635 ;
        RECT  3.955 1.905 4.115 3.105 ;
        RECT  1.545 2.945 3.955 3.105 ;
        RECT  3.615 0.585 3.775 1.295 ;
        RECT  3.615 1.870 3.775 2.765 ;
        RECT  2.975 0.585 3.615 0.745 ;
        RECT  2.455 2.605 3.615 2.765 ;
        RECT  3.275 1.095 3.435 2.425 ;
        RECT  3.155 1.095 3.275 1.255 ;
        RECT  2.825 2.265 3.275 2.425 ;
        RECT  2.895 0.925 3.155 1.255 ;
        RECT  2.815 0.495 2.975 0.745 ;
        RECT  1.750 0.925 2.895 1.085 ;
        RECT  2.465 0.495 2.815 0.655 ;
        RECT  2.455 1.265 2.595 2.215 ;
        RECT  2.435 1.265 2.455 2.765 ;
        RECT  2.325 1.265 2.435 1.425 ;
        RECT  2.295 2.055 2.435 2.765 ;
        RECT  2.195 2.055 2.295 2.585 ;
        RECT  1.995 1.615 2.255 1.875 ;
        RECT  1.775 2.055 2.195 2.215 ;
        RECT  1.410 1.615 1.995 1.775 ;
        RECT  1.515 1.955 1.775 2.215 ;
        RECT  1.590 0.460 1.750 1.085 ;
        RECT  1.135 0.460 1.590 0.620 ;
        RECT  1.385 2.425 1.545 3.105 ;
        RECT  1.250 0.830 1.410 1.775 ;
        RECT  1.295 2.425 1.385 2.585 ;
        RECT  1.135 1.955 1.295 2.585 ;
        RECT  0.525 0.830 1.250 0.990 ;
        RECT  0.945 2.845 1.205 3.105 ;
        RECT  1.070 1.955 1.135 2.215 ;
        RECT  1.035 1.200 1.070 2.215 ;
        RECT  0.910 1.200 1.035 2.125 ;
        RECT  0.725 2.845 0.945 3.005 ;
        RECT  0.735 1.200 0.910 1.360 ;
        RECT  0.565 1.615 0.725 3.005 ;
        RECT  0.525 1.615 0.565 1.775 ;
        RECT  0.365 0.830 0.525 1.775 ;
    END
END DFFXL

MACRO CMPR42X4
    CLASS CORE ;
    FOREIGN CMPR42X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  25.910 1.105 26.070 2.115 ;
        RECT  25.560 1.105 25.910 1.295 ;
        RECT  25.635 1.955 25.910 2.115 ;
        RECT  25.560 1.955 25.635 2.810 ;
        RECT  25.300 0.695 25.560 1.295 ;
        RECT  25.300 1.955 25.560 2.895 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.745 0.695 0.930 1.295 ;
        RECT  0.745 1.955 0.930 2.895 ;
        RECT  0.670 0.695 0.745 2.895 ;
        RECT  0.585 1.105 0.670 2.810 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.285 1.605 21.635 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.515 1.355 15.565 1.665 ;
        RECT  15.405 1.290 15.515 1.665 ;
        RECT  15.305 1.290 15.405 1.650 ;
        RECT  14.565 1.490 15.305 1.650 ;
        RECT  14.405 1.300 14.565 1.650 ;
        RECT  14.005 1.490 14.405 1.650 ;
        RECT  13.845 1.490 14.005 1.865 ;
        RECT  13.825 1.705 13.845 1.865 ;
        RECT  13.565 1.705 13.825 1.965 ;
        END
        ANTENNAGATEAREA     0.5083 ;
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.655 1.035 19.815 1.295 ;
        RECT  19.630 1.035 19.655 1.990 ;
        RECT  19.370 1.035 19.630 2.215 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.600 3.060 15.355 3.220 ;
        RECT  13.440 2.945 13.600 3.220 ;
        RECT  12.160 2.945 13.440 3.105 ;
        RECT  12.000 2.945 12.160 3.195 ;
        RECT  10.915 3.035 12.000 3.195 ;
        RECT  10.705 2.930 10.915 3.220 ;
        RECT  4.290 2.945 10.705 3.105 ;
        RECT  4.050 2.945 4.290 3.260 ;
        RECT  4.000 3.100 4.050 3.260 ;
        END
        ANTENNAGATEAREA     0.6786 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.580 1.705 9.840 2.055 ;
        RECT  8.615 1.895 9.580 2.055 ;
        RECT  8.540 1.895 8.615 2.175 ;
        RECT  8.380 1.895 8.540 2.765 ;
        RECT  7.090 2.605 8.380 2.765 ;
        RECT  6.930 1.895 7.090 2.765 ;
        RECT  2.175 1.895 6.930 2.055 ;
        RECT  2.150 1.700 2.175 2.055 ;
        RECT  1.990 1.695 2.150 2.055 ;
        RECT  1.965 1.695 1.990 1.990 ;
        RECT  1.890 1.695 1.965 1.955 ;
        END
        ANTENNAGATEAREA     1.2051 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.700 1.555 7.860 2.025 ;
        RECT  5.395 1.555 7.700 1.715 ;
        RECT  5.210 1.290 5.395 1.715 ;
        RECT  5.185 1.290 5.210 1.660 ;
        RECT  3.140 1.500 5.185 1.660 ;
        RECT  2.980 1.215 3.140 1.660 ;
        RECT  2.880 1.215 2.980 1.475 ;
        RECT  1.840 1.275 2.880 1.435 ;
        RECT  1.580 1.265 1.840 1.435 ;
        END
        ANTENNAGATEAREA     1.1037 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.070 -0.250 26.220 0.250 ;
        RECT  25.810 -0.250 26.070 0.830 ;
        RECT  25.020 -0.250 25.810 0.250 ;
        RECT  24.760 -0.250 25.020 0.405 ;
        RECT  23.320 -0.250 24.760 0.250 ;
        RECT  23.060 -0.250 23.320 0.405 ;
        RECT  21.360 -0.250 23.060 0.250 ;
        RECT  21.100 -0.250 21.360 0.405 ;
        RECT  20.355 -0.250 21.100 0.250 ;
        RECT  20.095 -0.250 20.355 0.405 ;
        RECT  19.275 -0.250 20.095 0.250 ;
        RECT  19.015 -0.250 19.275 0.405 ;
        RECT  15.415 -0.250 19.015 0.250 ;
        RECT  15.155 -0.250 15.415 0.405 ;
        RECT  12.645 -0.250 15.155 0.250 ;
        RECT  12.385 -0.250 12.645 0.405 ;
        RECT  10.380 -0.250 12.385 0.250 ;
        RECT  9.780 -0.250 10.380 0.405 ;
        RECT  8.130 -0.250 9.780 0.250 ;
        RECT  7.870 -0.250 8.130 0.865 ;
        RECT  7.260 -0.250 7.870 0.250 ;
        RECT  7.000 -0.250 7.260 1.375 ;
        RECT  6.210 -0.250 7.000 0.250 ;
        RECT  5.950 -0.250 6.210 0.405 ;
        RECT  5.120 -0.250 5.950 0.250 ;
        RECT  4.860 -0.250 5.120 0.405 ;
        RECT  3.340 -0.250 4.860 0.250 ;
        RECT  3.080 -0.250 3.340 0.405 ;
        RECT  1.470 -0.250 3.080 0.250 ;
        RECT  1.210 -0.250 1.470 0.745 ;
        RECT  0.390 -0.250 1.210 0.250 ;
        RECT  0.130 -0.250 0.390 1.295 ;
        RECT  0.000 -0.250 0.130 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.075 3.440 26.220 3.940 ;
        RECT  25.815 2.305 26.075 3.940 ;
        RECT  25.020 3.440 25.815 3.940 ;
        RECT  24.760 2.815 25.020 3.940 ;
        RECT  23.320 3.440 24.760 3.940 ;
        RECT  23.060 3.285 23.320 3.940 ;
        RECT  21.150 3.440 23.060 3.940 ;
        RECT  20.890 3.285 21.150 3.940 ;
        RECT  20.175 3.440 20.890 3.940 ;
        RECT  19.915 3.285 20.175 3.940 ;
        RECT  19.090 3.440 19.915 3.940 ;
        RECT  18.830 3.285 19.090 3.940 ;
        RECT  15.695 3.440 18.830 3.940 ;
        RECT  15.535 2.685 15.695 3.940 ;
        RECT  15.520 2.685 15.535 2.845 ;
        RECT  13.145 3.440 15.535 3.940 ;
        RECT  14.920 2.185 15.520 2.845 ;
        RECT  12.885 3.285 13.145 3.940 ;
        RECT  10.520 3.440 12.885 3.940 ;
        RECT  10.260 3.285 10.520 3.940 ;
        RECT  8.595 3.440 10.260 3.940 ;
        RECT  8.335 3.285 8.595 3.940 ;
        RECT  7.290 3.440 8.335 3.940 ;
        RECT  7.030 3.285 7.290 3.940 ;
        RECT  6.210 3.440 7.030 3.940 ;
        RECT  5.950 3.285 6.210 3.940 ;
        RECT  5.115 3.440 5.950 3.940 ;
        RECT  4.855 3.285 5.115 3.940 ;
        RECT  3.220 3.440 4.855 3.940 ;
        RECT  2.960 3.285 3.220 3.940 ;
        RECT  1.470 3.440 2.960 3.940 ;
        RECT  1.210 2.575 1.470 3.940 ;
        RECT  0.390 3.440 1.210 3.940 ;
        RECT  0.130 2.175 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  25.115 1.490 25.730 1.750 ;
        RECT  24.955 0.585 25.115 2.635 ;
        RECT  22.150 0.585 24.955 0.745 ;
        RECT  24.170 2.475 24.955 2.635 ;
        RECT  24.610 0.925 24.770 2.295 ;
        RECT  21.900 0.925 24.610 1.085 ;
        RECT  23.520 2.135 24.610 2.295 ;
        RECT  22.075 1.265 24.340 1.425 ;
        RECT  24.070 2.475 24.170 2.735 ;
        RECT  23.910 2.475 24.070 3.105 ;
        RECT  23.740 1.605 24.000 1.955 ;
        RECT  21.995 2.945 23.910 3.105 ;
        RECT  22.480 1.605 23.740 1.765 ;
        RECT  23.420 1.975 23.520 2.295 ;
        RECT  23.260 1.975 23.420 2.715 ;
        RECT  21.690 2.555 23.260 2.715 ;
        RECT  22.320 1.605 22.480 2.375 ;
        RECT  20.610 2.215 22.320 2.375 ;
        RECT  21.815 1.265 22.075 2.035 ;
        RECT  21.640 0.825 21.900 1.085 ;
        RECT  21.105 1.265 21.815 1.425 ;
        RECT  21.430 2.555 21.690 3.155 ;
        RECT  18.580 2.740 21.430 2.900 ;
        RECT  20.955 0.585 21.105 1.690 ;
        RECT  20.945 0.585 20.955 1.740 ;
        RECT  18.835 0.585 20.945 0.745 ;
        RECT  20.695 1.480 20.945 1.740 ;
        RECT  20.575 1.035 20.735 1.300 ;
        RECT  20.510 1.955 20.610 2.555 ;
        RECT  20.510 1.140 20.575 1.300 ;
        RECT  20.350 1.140 20.510 2.555 ;
        RECT  18.920 2.395 20.350 2.555 ;
        RECT  18.760 2.055 18.920 2.555 ;
        RECT  18.645 0.470 18.835 0.745 ;
        RECT  18.590 2.055 18.760 2.315 ;
        RECT  16.245 0.470 18.645 0.630 ;
        RECT  18.465 0.925 18.625 1.085 ;
        RECT  18.410 2.525 18.580 3.165 ;
        RECT  18.305 0.810 18.465 1.085 ;
        RECT  18.320 1.265 18.410 3.165 ;
        RECT  18.250 1.265 18.320 2.685 ;
        RECT  17.300 3.005 18.320 3.165 ;
        RECT  17.580 0.810 18.305 0.970 ;
        RECT  18.095 1.265 18.250 1.425 ;
        RECT  17.935 1.150 18.095 1.425 ;
        RECT  17.970 2.265 18.070 2.825 ;
        RECT  17.970 1.625 18.020 1.785 ;
        RECT  17.810 1.625 17.970 2.825 ;
        RECT  17.825 1.150 17.935 1.310 ;
        RECT  17.580 1.625 17.810 1.785 ;
        RECT  16.645 2.655 17.810 2.815 ;
        RECT  17.420 0.810 17.580 1.785 ;
        RECT  16.585 0.810 17.420 0.970 ;
        RECT  16.915 1.385 17.175 2.475 ;
        RECT  16.895 2.275 16.915 2.475 ;
        RECT  16.135 2.275 16.895 2.435 ;
        RECT  16.385 2.615 16.645 3.215 ;
        RECT  16.425 0.810 16.585 1.105 ;
        RECT  16.245 1.835 16.475 2.095 ;
        RECT  16.215 0.470 16.245 2.095 ;
        RECT  16.085 0.470 16.215 2.045 ;
        RECT  15.905 2.275 16.135 2.895 ;
        RECT  14.735 0.585 16.085 0.745 ;
        RECT  15.875 1.020 15.905 2.895 ;
        RECT  15.745 1.020 15.875 2.500 ;
        RECT  15.170 1.845 15.745 2.005 ;
        RECT  15.010 1.830 15.170 2.005 ;
        RECT  14.185 1.830 15.010 1.990 ;
        RECT  14.215 0.925 14.785 1.085 ;
        RECT  14.575 0.470 14.735 0.745 ;
        RECT  12.985 0.470 14.575 0.630 ;
        RECT  14.315 2.175 14.575 2.775 ;
        RECT  13.345 2.175 14.315 2.335 ;
        RECT  14.055 0.925 14.215 1.310 ;
        RECT  13.665 1.150 14.055 1.310 ;
        RECT  13.795 2.540 14.055 2.800 ;
        RECT  13.325 0.810 13.875 0.970 ;
        RECT  12.655 2.540 13.795 2.700 ;
        RECT  13.505 1.150 13.665 1.425 ;
        RECT  13.345 1.265 13.505 1.425 ;
        RECT  13.185 1.265 13.345 2.335 ;
        RECT  13.165 0.810 13.325 1.085 ;
        RECT  13.085 1.705 13.185 1.965 ;
        RECT  12.930 0.925 13.165 1.085 ;
        RECT  12.825 0.470 12.985 0.745 ;
        RECT  12.770 0.925 12.930 1.370 ;
        RECT  12.540 0.585 12.825 0.745 ;
        RECT  12.655 1.210 12.770 1.370 ;
        RECT  12.495 1.210 12.655 2.700 ;
        RECT  12.380 0.585 12.540 1.030 ;
        RECT  11.770 1.210 12.495 1.370 ;
        RECT  12.445 2.295 12.495 2.700 ;
        RECT  11.430 0.870 12.380 1.030 ;
        RECT  12.265 1.715 12.315 1.975 ;
        RECT  12.105 1.715 12.265 2.765 ;
        RECT  12.040 0.430 12.200 0.690 ;
        RECT  12.055 1.715 12.105 1.975 ;
        RECT  11.465 2.605 12.105 2.765 ;
        RECT  11.090 0.530 12.040 0.690 ;
        RECT  11.765 2.165 11.925 2.425 ;
        RECT  11.610 1.210 11.770 1.985 ;
        RECT  11.430 2.165 11.765 2.325 ;
        RECT  11.415 2.605 11.465 2.855 ;
        RECT  11.270 0.870 11.430 2.325 ;
        RECT  11.205 2.590 11.415 2.855 ;
        RECT  10.615 2.590 11.205 2.750 ;
        RECT  10.930 0.530 11.090 2.345 ;
        RECT  10.710 0.530 10.930 0.790 ;
        RECT  10.800 2.185 10.930 2.345 ;
        RECT  10.615 1.010 10.750 2.000 ;
        RECT  10.590 1.010 10.615 2.750 ;
        RECT  10.525 1.010 10.590 1.170 ;
        RECT  10.455 1.840 10.590 2.750 ;
        RECT  10.365 0.875 10.525 1.170 ;
        RECT  9.410 2.590 10.455 2.750 ;
        RECT  9.190 0.875 10.365 1.035 ;
        RECT  10.180 1.400 10.320 1.660 ;
        RECT  10.020 1.215 10.180 2.400 ;
        RECT  8.680 1.215 10.020 1.375 ;
        RECT  9.160 2.240 10.020 2.400 ;
        RECT  8.200 1.555 9.330 1.715 ;
        RECT  8.930 0.775 9.190 1.035 ;
        RECT  8.900 2.240 9.160 2.500 ;
        RECT  8.520 0.685 8.680 1.375 ;
        RECT  8.420 0.685 8.520 0.945 ;
        RECT  8.040 1.165 8.200 2.425 ;
        RECT  7.510 1.165 8.040 1.325 ;
        RECT  7.510 2.265 8.040 2.425 ;
        RECT  6.490 0.765 6.750 1.365 ;
        RECT  6.490 2.235 6.750 2.765 ;
        RECT  5.620 0.785 6.490 1.045 ;
        RECT  5.670 2.235 6.490 2.495 ;
        RECT  5.410 2.235 5.670 2.765 ;
        RECT  5.410 0.755 5.620 1.045 ;
        RECT  3.990 0.755 5.410 0.915 ;
        RECT  3.830 2.235 5.410 2.395 ;
        RECT  3.710 1.095 4.760 1.255 ;
        RECT  3.580 2.575 4.600 2.735 ;
        RECT  3.450 0.705 3.710 1.305 ;
        RECT  3.320 2.390 3.580 2.735 ;
        RECT  2.490 0.705 3.450 0.865 ;
        RECT  2.360 2.575 3.320 2.735 ;
        RECT  2.230 0.495 2.490 1.095 ;
        RECT  2.100 2.235 2.360 2.835 ;
        RECT  1.400 0.925 2.230 1.085 ;
        RECT  1.400 2.235 2.100 2.395 ;
        RECT  1.240 0.925 1.400 2.395 ;
        RECT  0.925 1.480 1.240 1.740 ;
    END
END CMPR42X4

MACRO CMPR42X2
    CLASS CORE ;
    FOREIGN CMPR42X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.270 0.695 18.275 1.295 ;
        RECT  18.270 2.110 18.275 2.895 ;
        RECT  18.110 0.695 18.270 2.895 ;
        RECT  18.015 0.695 18.110 1.295 ;
        RECT  18.010 1.955 18.110 2.895 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 0.695 0.520 1.295 ;
        RECT  0.335 1.920 0.390 2.895 ;
        RECT  0.260 0.695 0.335 2.895 ;
        RECT  0.125 1.105 0.260 2.895 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.515 1.585 15.700 1.945 ;
        RECT  15.305 1.585 15.515 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.835 1.355 11.870 1.665 ;
        RECT  11.710 1.290 11.835 1.665 ;
        RECT  11.625 1.290 11.710 1.650 ;
        RECT  10.870 1.490 11.625 1.650 ;
        RECT  10.710 1.300 10.870 1.650 ;
        RECT  10.310 1.490 10.710 1.650 ;
        RECT  10.150 1.490 10.310 1.865 ;
        RECT  10.130 1.705 10.150 1.865 ;
        RECT  9.870 1.705 10.130 1.965 ;
        END
        ANTENNAGATEAREA     0.5044 ;
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.145 1.035 14.180 1.295 ;
        RECT  13.920 1.035 14.145 2.215 ;
        END
        ANTENNADIFFAREA     0.5794 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.840 3.060 11.660 3.220 ;
        RECT  9.680 2.945 9.840 3.220 ;
        RECT  8.730 2.945 9.680 3.105 ;
        RECT  8.570 2.945 8.730 3.195 ;
        RECT  7.235 3.035 8.570 3.195 ;
        RECT  7.025 2.930 7.235 3.220 ;
        RECT  7.010 2.945 7.025 3.220 ;
        RECT  2.210 2.945 7.010 3.105 ;
        RECT  2.000 2.945 2.210 3.260 ;
        RECT  1.950 3.100 2.000 3.260 ;
        END
        ANTENNAGATEAREA     0.4654 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.100 1.705 6.150 1.965 ;
        RECT  5.890 1.705 6.100 2.055 ;
        RECT  5.000 1.895 5.890 2.055 ;
        RECT  4.840 1.895 5.000 2.765 ;
        RECT  3.770 2.605 4.840 2.765 ;
        RECT  3.610 1.895 3.770 2.765 ;
        RECT  1.715 1.895 3.610 2.055 ;
        RECT  1.610 1.700 1.715 2.055 ;
        RECT  1.530 1.695 1.610 2.055 ;
        RECT  1.505 1.695 1.530 1.990 ;
        RECT  1.350 1.695 1.505 1.955 ;
        END
        ANTENNAGATEAREA     0.7787 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 1.555 4.320 2.075 ;
        RECT  2.805 1.555 4.160 1.715 ;
        RECT  2.635 1.355 2.805 1.715 ;
        RECT  2.610 1.290 2.635 1.715 ;
        RECT  2.540 1.280 2.610 1.715 ;
        RECT  2.425 1.280 2.540 1.580 ;
        RECT  1.300 1.280 2.425 1.440 ;
        RECT  1.040 1.265 1.300 1.440 ;
        END
        ANTENNAGATEAREA     0.6773 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.735 -0.250 18.400 0.250 ;
        RECT  17.475 -0.250 17.735 0.405 ;
        RECT  15.835 -0.250 17.475 0.250 ;
        RECT  15.575 -0.250 15.835 0.405 ;
        RECT  14.720 -0.250 15.575 0.250 ;
        RECT  14.460 -0.250 14.720 0.405 ;
        RECT  11.775 -0.250 14.460 0.250 ;
        RECT  11.515 -0.250 11.775 0.405 ;
        RECT  8.950 -0.250 11.515 0.250 ;
        RECT  8.690 -0.250 8.950 0.405 ;
        RECT  6.720 -0.250 8.690 0.250 ;
        RECT  6.520 -0.250 6.720 0.795 ;
        RECT  6.120 -0.250 6.520 0.405 ;
        RECT  4.480 -0.250 6.120 0.250 ;
        RECT  4.220 -0.250 4.480 0.945 ;
        RECT  3.000 -0.250 4.220 0.250 ;
        RECT  2.740 -0.250 3.000 0.745 ;
        RECT  1.060 -0.250 2.740 0.250 ;
        RECT  0.800 -0.250 1.060 0.745 ;
        RECT  0.000 -0.250 0.800 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.690 3.440 18.400 3.940 ;
        RECT  17.430 3.285 17.690 3.940 ;
        RECT  15.465 3.440 17.430 3.940 ;
        RECT  14.425 3.285 15.465 3.940 ;
        RECT  12.000 3.440 14.425 3.940 ;
        RECT  11.840 2.685 12.000 3.940 ;
        RECT  11.825 2.685 11.840 2.845 ;
        RECT  9.320 3.440 11.840 3.940 ;
        RECT  11.225 2.185 11.825 2.845 ;
        RECT  9.060 3.285 9.320 3.940 ;
        RECT  6.830 3.440 9.060 3.940 ;
        RECT  6.570 3.285 6.830 3.940 ;
        RECT  4.850 3.440 6.570 3.940 ;
        RECT  4.590 3.285 4.850 3.940 ;
        RECT  3.840 3.440 4.590 3.940 ;
        RECT  3.580 3.285 3.840 3.940 ;
        RECT  2.750 3.440 3.580 3.940 ;
        RECT  2.490 3.285 2.750 3.940 ;
        RECT  0.930 3.440 2.490 3.940 ;
        RECT  0.670 2.575 0.930 3.940 ;
        RECT  0.000 3.440 0.670 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.830 1.500 17.920 1.760 ;
        RECT  17.670 0.585 17.830 2.965 ;
        RECT  16.625 0.585 17.670 0.745 ;
        RECT  16.410 2.805 17.670 2.965 ;
        RECT  17.235 0.925 17.395 1.955 ;
        RECT  16.425 0.925 17.235 1.085 ;
        RECT  17.220 1.695 17.235 1.955 ;
        RECT  17.060 1.695 17.220 2.625 ;
        RECT  16.230 2.465 17.060 2.625 ;
        RECT  16.265 1.265 17.055 1.425 ;
        RECT  16.645 1.745 16.745 2.005 ;
        RECT  16.485 1.745 16.645 2.285 ;
        RECT  15.890 2.125 16.485 2.285 ;
        RECT  16.265 0.805 16.425 1.085 ;
        RECT  16.115 0.805 16.265 1.065 ;
        RECT  16.085 1.265 16.265 1.935 ;
        RECT  16.070 2.465 16.230 2.715 ;
        RECT  16.005 1.245 16.085 1.935 ;
        RECT  16.040 2.555 16.070 2.715 ;
        RECT  15.780 2.555 16.040 3.155 ;
        RECT  15.925 1.245 16.005 1.520 ;
        RECT  15.835 1.245 15.925 1.405 ;
        RECT  15.730 2.125 15.890 2.330 ;
        RECT  15.675 0.585 15.835 1.405 ;
        RECT  13.530 2.895 15.780 3.055 ;
        RECT  15.120 2.170 15.730 2.330 ;
        RECT  14.780 0.585 15.675 0.745 ;
        RECT  15.120 1.035 15.260 1.295 ;
        RECT  14.960 1.035 15.120 2.555 ;
        RECT  14.835 2.265 14.960 2.555 ;
        RECT  13.885 2.395 14.835 2.555 ;
        RECT  14.620 0.585 14.780 1.665 ;
        RECT  14.160 0.585 14.620 0.745 ;
        RECT  14.000 0.470 14.160 0.745 ;
        RECT  12.660 0.470 14.000 0.630 ;
        RECT  13.625 2.395 13.885 2.655 ;
        RECT  13.580 0.945 13.740 2.170 ;
        RECT  13.560 0.945 13.580 1.105 ;
        RECT  13.430 2.010 13.580 2.170 ;
        RECT  13.300 0.845 13.560 1.105 ;
        RECT  13.430 2.895 13.530 3.155 ;
        RECT  13.270 2.010 13.430 3.155 ;
        RECT  13.010 1.535 13.400 1.795 ;
        RECT  13.000 1.535 13.010 3.070 ;
        RECT  12.840 0.845 13.000 3.070 ;
        RECT  12.750 2.470 12.840 3.070 ;
        RECT  12.550 0.470 12.660 1.915 ;
        RECT  12.500 0.470 12.550 2.015 ;
        RECT  10.595 0.585 12.500 0.745 ;
        RECT  12.390 1.755 12.500 2.015 ;
        RECT  12.210 2.345 12.440 3.070 ;
        RECT  12.210 1.020 12.320 1.280 ;
        RECT  12.180 1.020 12.210 3.070 ;
        RECT  12.050 1.020 12.180 2.505 ;
        RECT  11.475 1.845 12.050 2.005 ;
        RECT  11.315 1.830 11.475 2.005 ;
        RECT  10.490 1.830 11.315 1.990 ;
        RECT  10.520 0.925 11.090 1.085 ;
        RECT  10.620 2.175 10.880 2.775 ;
        RECT  9.650 2.175 10.620 2.335 ;
        RECT  10.435 0.470 10.595 0.745 ;
        RECT  10.360 0.925 10.520 1.310 ;
        RECT  9.290 0.470 10.435 0.630 ;
        RECT  9.970 1.150 10.360 1.310 ;
        RECT  10.100 2.540 10.360 2.800 ;
        RECT  9.630 0.810 10.180 0.970 ;
        RECT  8.960 2.540 10.100 2.700 ;
        RECT  9.810 1.150 9.970 1.425 ;
        RECT  9.650 1.265 9.810 1.425 ;
        RECT  9.490 1.265 9.650 2.335 ;
        RECT  9.470 0.810 9.630 1.085 ;
        RECT  9.390 1.705 9.490 1.965 ;
        RECT  9.195 0.925 9.470 1.085 ;
        RECT  9.130 0.470 9.290 0.745 ;
        RECT  9.035 0.925 9.195 1.370 ;
        RECT  8.850 0.585 9.130 0.745 ;
        RECT  8.960 1.210 9.035 1.370 ;
        RECT  8.800 1.210 8.960 2.700 ;
        RECT  8.690 0.585 8.850 1.030 ;
        RECT  8.080 1.210 8.800 1.370 ;
        RECT  8.750 2.295 8.800 2.700 ;
        RECT  7.740 0.870 8.690 1.030 ;
        RECT  8.570 1.715 8.620 1.975 ;
        RECT  8.410 1.715 8.570 2.765 ;
        RECT  8.350 0.430 8.510 0.690 ;
        RECT  8.360 1.715 8.410 1.975 ;
        RECT  7.770 2.605 8.410 2.765 ;
        RECT  7.400 0.530 8.350 0.690 ;
        RECT  8.070 2.165 8.230 2.425 ;
        RECT  7.920 1.210 8.080 1.985 ;
        RECT  7.740 2.165 8.070 2.325 ;
        RECT  7.720 2.605 7.770 2.855 ;
        RECT  7.580 0.870 7.740 2.325 ;
        RECT  7.510 2.590 7.720 2.855 ;
        RECT  6.870 2.590 7.510 2.750 ;
        RECT  7.240 0.530 7.400 2.345 ;
        RECT  7.020 0.570 7.240 0.830 ;
        RECT  7.110 2.185 7.240 2.345 ;
        RECT  6.900 1.010 7.060 2.005 ;
        RECT  6.340 1.010 6.900 1.170 ;
        RECT  6.870 1.845 6.900 2.005 ;
        RECT  6.710 1.845 6.870 2.750 ;
        RECT  5.720 2.590 6.710 2.750 ;
        RECT  6.530 1.405 6.630 1.665 ;
        RECT  6.370 1.355 6.530 2.400 ;
        RECT  6.000 1.355 6.370 1.515 ;
        RECT  5.470 2.240 6.370 2.400 ;
        RECT  6.180 0.875 6.340 1.170 ;
        RECT  5.500 0.875 6.180 1.035 ;
        RECT  5.840 1.215 6.000 1.515 ;
        RECT  5.000 1.215 5.840 1.375 ;
        RECT  4.660 1.555 5.660 1.715 ;
        RECT  5.240 0.775 5.500 1.035 ;
        RECT  5.210 2.240 5.470 2.760 ;
        RECT  4.840 0.685 5.000 1.375 ;
        RECT  4.730 0.685 4.840 0.945 ;
        RECT  4.500 1.215 4.660 2.425 ;
        RECT  3.940 1.215 4.500 1.375 ;
        RECT  4.000 2.265 4.500 2.425 ;
        RECT  3.680 1.115 3.940 1.375 ;
        RECT  3.440 0.605 3.540 0.865 ;
        RECT  3.280 0.605 3.440 1.095 ;
        RECT  3.030 2.265 3.290 2.765 ;
        RECT  2.460 0.935 3.280 1.095 ;
        RECT  2.380 2.265 3.030 2.425 ;
        RECT  2.200 0.495 2.460 1.095 ;
        RECT  2.120 2.265 2.380 2.595 ;
        RECT  1.690 0.495 1.950 1.095 ;
        RECT  1.560 2.235 1.820 2.835 ;
        RECT  0.860 0.925 1.690 1.085 ;
        RECT  0.860 2.235 1.560 2.395 ;
        RECT  0.700 0.925 0.860 2.395 ;
        RECT  0.560 1.480 0.700 1.740 ;
    END
END CMPR42X2

MACRO CMPR42X1
    CLASS CORE ;
    FOREIGN CMPR42X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.560 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.435 1.035 16.440 2.335 ;
        RECT  16.430 1.035 16.435 2.400 ;
        RECT  16.280 1.035 16.430 2.555 ;
        RECT  16.170 1.035 16.280 1.295 ;
        RECT  16.170 1.955 16.280 2.555 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 0.795 0.680 1.055 ;
        RECT  0.420 0.795 0.580 1.300 ;
        RECT  0.285 1.140 0.420 1.300 ;
        RECT  0.285 1.955 0.390 2.555 ;
        RECT  0.130 1.140 0.285 2.555 ;
        RECT  0.125 1.140 0.130 2.400 ;
        END
        ANTENNADIFFAREA     0.3646 ;
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.925 2.425 14.135 2.810 ;
        RECT  13.630 2.425 13.925 2.635 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.545 1.355 10.550 1.650 ;
        RECT  10.455 1.300 10.545 1.650 ;
        RECT  10.245 1.290 10.455 1.650 ;
        RECT  10.185 1.300 10.245 1.650 ;
        END
        ANTENNAGATEAREA     0.3484 ;
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.950 1.290 13.215 1.580 ;
        RECT  12.800 1.100 12.950 1.580 ;
        RECT  12.690 1.100 12.800 2.295 ;
        RECT  12.540 1.290 12.690 2.295 ;
        END
        ANTENNADIFFAREA     0.3230 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.920 3.005 10.120 3.165 ;
        RECT  8.760 2.940 8.920 3.165 ;
        RECT  7.695 2.940 8.760 3.100 ;
        RECT  7.485 2.930 7.695 3.220 ;
        RECT  6.735 3.050 7.485 3.210 ;
        RECT  6.575 2.945 6.735 3.210 ;
        RECT  1.990 2.945 6.575 3.105 ;
        RECT  1.730 2.895 1.990 3.155 ;
        END
        ANTENNAGATEAREA     0.2795 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.330 1.770 5.590 2.055 ;
        RECT  4.545 1.895 5.330 2.055 ;
        RECT  4.385 1.895 4.545 2.765 ;
        RECT  3.380 2.605 4.385 2.765 ;
        RECT  3.280 1.990 3.380 2.765 ;
        RECT  3.220 1.865 3.280 2.765 ;
        RECT  3.120 1.865 3.220 2.250 ;
        RECT  1.715 1.865 3.120 2.025 ;
        RECT  1.505 1.700 1.715 2.025 ;
        RECT  1.485 1.865 1.505 2.025 ;
        RECT  1.225 1.865 1.485 2.125 ;
        END
        ANTENNAGATEAREA     0.4407 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.700 1.525 3.860 1.965 ;
        RECT  3.095 1.525 3.700 1.685 ;
        RECT  2.960 1.515 3.095 1.685 ;
        RECT  2.750 1.285 2.960 1.685 ;
        RECT  2.700 1.285 2.750 1.580 ;
        RECT  2.425 1.290 2.700 1.580 ;
        RECT  1.460 1.290 2.425 1.450 ;
        RECT  1.250 1.280 1.460 1.450 ;
        RECT  1.200 1.280 1.250 1.440 ;
        END
        ANTENNAGATEAREA     0.3848 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.030 -0.250 16.560 0.250 ;
        RECT  15.770 -0.250 16.030 0.405 ;
        RECT  13.840 -0.250 15.770 0.250 ;
        RECT  13.240 -0.250 13.840 0.405 ;
        RECT  10.515 -0.250 13.240 0.250 ;
        RECT  10.355 -0.250 10.515 0.770 ;
        RECT  8.510 -0.250 10.355 0.250 ;
        RECT  8.250 -0.250 8.510 0.405 ;
        RECT  6.090 -0.250 8.250 0.250 ;
        RECT  5.830 -0.250 6.090 0.405 ;
        RECT  4.300 -0.250 5.830 0.250 ;
        RECT  4.040 -0.250 4.300 0.945 ;
        RECT  3.160 -0.250 4.040 0.250 ;
        RECT  2.900 -0.250 3.160 0.405 ;
        RECT  1.260 -0.250 2.900 0.250 ;
        RECT  1.000 -0.250 1.260 0.745 ;
        RECT  0.000 -0.250 1.000 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.030 3.440 16.560 3.940 ;
        RECT  15.770 3.285 16.030 3.940 ;
        RECT  13.350 3.440 15.770 3.940 ;
        RECT  13.090 3.285 13.350 3.940 ;
        RECT  10.490 3.440 13.090 3.940 ;
        RECT  10.330 2.225 10.490 3.940 ;
        RECT  10.230 2.225 10.330 2.825 ;
        RECT  8.580 3.440 10.330 3.940 ;
        RECT  8.320 3.285 8.580 3.940 ;
        RECT  6.250 3.440 8.320 3.940 ;
        RECT  5.990 3.285 6.250 3.940 ;
        RECT  4.380 3.440 5.990 3.940 ;
        RECT  4.120 3.285 4.380 3.940 ;
        RECT  3.590 3.440 4.120 3.940 ;
        RECT  3.330 3.285 3.590 3.940 ;
        RECT  2.460 3.440 3.330 3.940 ;
        RECT  2.200 3.285 2.460 3.940 ;
        RECT  0.790 3.440 2.200 3.940 ;
        RECT  0.530 2.875 0.790 3.940 ;
        RECT  0.000 3.440 0.530 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.990 1.500 16.080 1.760 ;
        RECT  15.830 0.585 15.990 3.055 ;
        RECT  14.910 0.585 15.830 0.745 ;
        RECT  15.170 2.895 15.830 3.055 ;
        RECT  15.440 0.925 15.600 2.670 ;
        RECT  14.660 0.925 15.440 1.085 ;
        RECT  14.660 2.510 15.440 2.670 ;
        RECT  15.100 1.265 15.260 2.330 ;
        RECT  14.910 2.895 15.170 3.155 ;
        RECT  14.070 1.265 15.100 1.425 ;
        RECT  13.445 2.085 15.100 2.245 ;
        RECT  13.730 1.745 14.830 1.905 ;
        RECT  14.500 0.525 14.660 1.085 ;
        RECT  14.560 2.510 14.660 2.985 ;
        RECT  14.500 2.510 14.560 3.150 ;
        RECT  14.400 0.525 14.500 0.785 ;
        RECT  14.400 2.725 14.500 3.150 ;
        RECT  13.735 2.990 14.400 3.150 ;
        RECT  13.910 1.115 14.070 1.425 ;
        RECT  13.575 2.945 13.735 3.150 ;
        RECT  13.570 0.585 13.730 1.905 ;
        RECT  12.905 2.945 13.575 3.105 ;
        RECT  12.780 0.585 13.570 0.745 ;
        RECT  13.285 2.085 13.445 2.765 ;
        RECT  12.560 2.605 13.285 2.765 ;
        RECT  12.745 2.945 12.905 3.210 ;
        RECT  12.620 0.470 12.780 0.745 ;
        RECT  12.100 3.050 12.745 3.210 ;
        RECT  11.540 0.470 12.620 0.630 ;
        RECT  12.400 2.605 12.560 2.820 ;
        RECT  12.360 0.850 12.440 1.010 ;
        RECT  12.280 2.660 12.400 2.820 ;
        RECT  12.220 0.850 12.360 2.130 ;
        RECT  12.200 0.850 12.220 2.480 ;
        RECT  12.180 0.850 12.200 1.010 ;
        RECT  12.100 1.970 12.200 2.480 ;
        RECT  12.060 1.970 12.100 3.210 ;
        RECT  11.940 2.320 12.060 3.210 ;
        RECT  11.880 1.500 12.020 1.760 ;
        RECT  11.720 0.810 11.880 2.140 ;
        RECT  11.630 1.980 11.720 2.140 ;
        RECT  11.470 1.980 11.630 2.515 ;
        RECT  11.380 0.470 11.540 1.800 ;
        RECT  11.370 2.255 11.470 2.515 ;
        RECT  10.855 0.680 11.380 0.840 ;
        RECT  11.230 1.640 11.380 1.800 ;
        RECT  11.070 1.640 11.230 1.970 ;
        RECT  11.040 1.020 11.200 1.460 ;
        RECT  10.890 2.250 11.110 2.510 ;
        RECT  10.890 1.300 11.040 1.460 ;
        RECT  10.850 1.300 10.890 2.510 ;
        RECT  10.695 0.680 10.855 1.110 ;
        RECT  10.730 1.300 10.850 2.410 ;
        RECT  9.780 1.835 10.730 1.995 ;
        RECT  10.170 0.950 10.695 1.110 ;
        RECT  10.010 0.505 10.170 1.110 ;
        RECT  9.135 0.505 10.010 0.665 ;
        RECT  9.690 2.175 9.950 2.775 ;
        RECT  9.670 0.850 9.830 1.500 ;
        RECT  9.520 1.705 9.780 1.995 ;
        RECT  9.340 2.175 9.690 2.335 ;
        RECT  9.340 1.340 9.670 1.500 ;
        RECT  9.180 2.545 9.440 2.805 ;
        RECT  8.220 0.925 9.370 1.085 ;
        RECT  9.180 1.340 9.340 2.335 ;
        RECT  8.460 1.635 9.180 1.895 ;
        RECT  8.220 2.590 9.180 2.750 ;
        RECT  8.975 0.505 9.135 0.745 ;
        RECT  7.640 0.585 8.975 0.745 ;
        RECT  8.060 0.925 8.220 2.750 ;
        RECT  7.890 1.020 8.060 1.280 ;
        RECT  7.960 1.710 8.060 2.750 ;
        RECT  7.360 1.710 7.960 1.970 ;
        RECT  7.450 2.150 7.710 2.750 ;
        RECT  7.540 0.585 7.640 1.145 ;
        RECT  7.480 0.585 7.540 1.460 ;
        RECT  7.380 0.885 7.480 1.460 ;
        RECT  7.180 2.150 7.450 2.310 ;
        RECT  7.180 1.300 7.380 1.460 ;
        RECT  6.940 2.605 7.200 2.870 ;
        RECT  7.020 1.300 7.180 2.310 ;
        RECT  6.840 0.835 7.130 1.095 ;
        RECT  6.410 2.605 6.940 2.765 ;
        RECT  6.680 0.530 6.840 2.405 ;
        RECT  6.430 0.530 6.680 0.690 ;
        RECT  6.590 2.145 6.680 2.405 ;
        RECT  6.410 1.635 6.500 1.895 ;
        RECT  6.270 0.430 6.430 0.690 ;
        RECT  6.250 0.870 6.410 2.765 ;
        RECT  5.120 0.870 6.250 1.030 ;
        RECT  5.230 2.605 6.250 2.765 ;
        RECT  5.970 1.420 6.070 2.425 ;
        RECT  5.910 1.215 5.970 2.425 ;
        RECT  5.810 1.215 5.910 1.680 ;
        RECT  4.885 2.265 5.910 2.425 ;
        RECT  4.840 1.215 5.810 1.375 ;
        RECT  4.205 1.555 5.105 1.715 ;
        RECT  4.725 2.265 4.885 2.525 ;
        RECT  4.680 0.770 4.840 1.375 ;
        RECT  4.580 0.770 4.680 1.030 ;
        RECT  4.045 1.125 4.205 2.425 ;
        RECT  3.730 1.125 4.045 1.285 ;
        RECT  3.760 2.265 4.045 2.425 ;
        RECT  3.470 1.025 3.730 1.285 ;
        RECT  3.440 0.515 3.700 0.775 ;
        RECT  2.620 0.615 3.440 0.775 ;
        RECT  2.935 2.600 3.040 2.760 ;
        RECT  2.775 2.335 2.935 2.760 ;
        RECT  2.190 2.335 2.775 2.495 ;
        RECT  2.460 0.615 2.620 1.045 ;
        RECT  2.360 0.785 2.460 1.045 ;
        RECT  1.930 2.235 2.190 2.495 ;
        RECT  1.850 0.785 2.110 1.095 ;
        RECT  1.020 0.935 1.850 1.095 ;
        RECT  1.390 2.330 1.650 2.590 ;
        RECT  1.020 2.330 1.390 2.490 ;
        RECT  0.860 0.935 1.020 2.490 ;
        RECT  0.480 1.480 0.860 1.740 ;
    END
END CMPR42X1

MACRO AHCSHCONX4
    CLASS CORE ;
    FOREIGN AHCSHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.145 2.110 8.155 2.810 ;
        RECT  8.105 0.915 8.145 2.810 ;
        RECT  7.985 0.695 8.105 2.940 ;
        RECT  7.845 0.695 7.985 1.295 ;
        RECT  7.845 2.000 7.985 2.940 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.995 2.405 7.395 2.810 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.240 1.815 2.895 ;
        RECT  1.255 2.240 1.505 2.400 ;
        RECT  1.255 0.850 1.305 1.110 ;
        RECT  1.045 0.850 1.255 2.400 ;
        RECT  0.795 2.240 1.045 2.400 ;
        RECT  0.525 2.240 0.795 2.895 ;
        END
        ANTENNADIFFAREA     1.2567 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.965 1.665 3.125 2.665 ;
        RECT  2.955 1.665 2.965 1.825 ;
        RECT  2.190 2.505 2.965 2.665 ;
        RECT  2.795 1.555 2.955 1.825 ;
        RECT  2.030 1.870 2.190 2.665 ;
        RECT  1.715 1.870 2.030 2.030 ;
        RECT  1.515 1.290 1.715 2.030 ;
        RECT  1.505 1.290 1.515 1.805 ;
        RECT  1.465 1.545 1.505 1.805 ;
        END
        ANTENNAGATEAREA     0.8242 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.055 1.290 2.235 1.690 ;
        RECT  1.895 0.950 2.055 1.690 ;
        RECT  1.840 0.950 1.895 1.110 ;
        RECT  1.680 0.510 1.840 1.110 ;
        RECT  0.865 0.510 1.680 0.670 ;
        RECT  0.705 0.510 0.865 1.565 ;
        RECT  0.645 1.405 0.705 1.565 ;
        RECT  0.385 1.405 0.645 1.665 ;
        END
        ANTENNAGATEAREA     0.7540 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.555 -0.250 8.280 0.250 ;
        RECT  7.295 -0.250 7.555 0.405 ;
        RECT  4.925 -0.250 7.295 0.250 ;
        RECT  4.665 -0.250 4.925 0.575 ;
        RECT  2.325 -0.250 4.665 0.250 ;
        RECT  2.065 -0.250 2.325 0.740 ;
        RECT  0.475 -0.250 2.065 0.250 ;
        RECT  0.215 -0.250 0.475 1.075 ;
        RECT  0.000 -0.250 0.215 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.555 3.440 8.280 3.940 ;
        RECT  7.295 3.285 7.555 3.940 ;
        RECT  4.795 3.440 7.295 3.940 ;
        RECT  4.535 3.115 4.795 3.940 ;
        RECT  2.325 3.440 4.535 3.940 ;
        RECT  2.065 2.955 2.325 3.940 ;
        RECT  1.295 3.440 2.065 3.940 ;
        RECT  1.035 2.615 1.295 3.940 ;
        RECT  0.385 3.440 1.035 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.545 1.525 7.805 1.785 ;
        RECT  7.465 1.525 7.545 1.685 ;
        RECT  7.305 0.695 7.465 1.685 ;
        RECT  6.955 0.695 7.305 0.855 ;
        RECT  7.025 1.955 7.155 2.215 ;
        RECT  7.025 1.035 7.125 1.295 ;
        RECT  6.865 1.035 7.025 2.215 ;
        RECT  6.795 0.495 6.955 0.855 ;
        RECT  6.630 1.525 6.865 1.785 ;
        RECT  6.105 0.495 6.795 0.655 ;
        RECT  6.445 0.835 6.615 1.095 ;
        RECT  6.445 2.065 6.615 3.005 ;
        RECT  6.285 0.835 6.445 3.160 ;
        RECT  5.135 3.000 6.285 3.160 ;
        RECT  5.945 0.495 6.105 2.645 ;
        RECT  5.845 0.495 5.945 1.095 ;
        RECT  5.845 2.045 5.945 2.645 ;
        RECT  5.435 0.475 5.595 2.815 ;
        RECT  5.335 0.475 5.435 0.915 ;
        RECT  5.335 2.555 5.435 2.815 ;
        RECT  4.485 0.755 5.335 0.915 ;
        RECT  5.095 1.095 5.195 2.305 ;
        RECT  4.975 2.775 5.135 3.160 ;
        RECT  5.035 1.095 5.095 2.595 ;
        RECT  4.935 1.095 5.035 1.255 ;
        RECT  4.935 2.045 5.035 2.595 ;
        RECT  3.465 2.775 4.975 2.935 ;
        RECT  3.805 2.435 4.935 2.595 ;
        RECT  4.325 0.625 4.485 1.690 ;
        RECT  2.935 0.625 4.325 0.785 ;
        RECT  4.145 2.095 4.245 2.255 ;
        RECT  3.985 0.985 4.145 2.255 ;
        RECT  3.645 1.675 3.805 2.595 ;
        RECT  3.465 0.965 3.660 1.225 ;
        RECT  3.305 0.965 3.465 2.985 ;
        RECT  2.675 0.625 2.935 1.245 ;
        RECT  2.625 2.005 2.785 2.295 ;
        RECT  2.615 1.085 2.675 1.245 ;
        RECT  2.615 2.005 2.625 2.165 ;
        RECT  2.455 1.085 2.615 2.165 ;
    END
END AHCSHCONX4

MACRO AHCSHCONX2
    CLASS CORE ;
    FOREIGN AHCSHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.225 0.695 7.235 1.105 ;
        RECT  7.225 2.110 7.235 2.940 ;
        RECT  7.065 0.695 7.225 2.940 ;
        RECT  6.925 0.695 7.065 1.295 ;
        RECT  6.925 2.000 7.065 2.940 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.075 2.405 6.475 2.810 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 2.240 0.895 2.895 ;
        RECT  0.335 2.240 0.585 2.400 ;
        RECT  0.320 0.475 0.580 1.075 ;
        RECT  0.285 2.110 0.335 2.400 ;
        RECT  0.285 0.915 0.320 1.075 ;
        RECT  0.125 0.915 0.285 2.400 ;
        END
        ANTENNADIFFAREA     0.6572 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 1.665 2.205 2.635 ;
        RECT  2.035 1.665 2.045 1.825 ;
        RECT  1.235 2.475 2.045 2.635 ;
        RECT  1.875 1.555 2.035 1.825 ;
        RECT  1.075 1.870 1.235 2.635 ;
        RECT  0.795 1.870 1.075 2.030 ;
        RECT  0.595 1.290 0.795 2.030 ;
        RECT  0.585 1.290 0.595 1.805 ;
        RECT  0.495 1.545 0.585 1.805 ;
        END
        ANTENNAGATEAREA     0.5876 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.975 1.290 1.315 1.690 ;
        END
        ANTENNAGATEAREA     0.5174 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.635 -0.250 7.360 0.250 ;
        RECT  6.375 -0.250 6.635 0.405 ;
        RECT  4.005 -0.250 6.375 0.250 ;
        RECT  3.745 -0.250 4.005 0.575 ;
        RECT  1.405 -0.250 3.745 0.250 ;
        RECT  1.145 -0.250 1.405 1.030 ;
        RECT  0.000 -0.250 1.145 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.635 3.440 7.360 3.940 ;
        RECT  6.375 3.285 6.635 3.940 ;
        RECT  3.875 3.440 6.375 3.940 ;
        RECT  3.615 3.115 3.875 3.940 ;
        RECT  1.405 3.440 3.615 3.940 ;
        RECT  1.145 2.865 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.615 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.625 1.525 6.885 1.785 ;
        RECT  6.545 1.525 6.625 1.685 ;
        RECT  6.385 0.695 6.545 1.685 ;
        RECT  6.035 0.695 6.385 0.855 ;
        RECT  6.105 1.955 6.235 2.215 ;
        RECT  6.105 1.035 6.205 1.295 ;
        RECT  5.945 1.035 6.105 2.215 ;
        RECT  5.875 0.495 6.035 0.855 ;
        RECT  5.710 1.525 5.945 1.785 ;
        RECT  5.185 0.495 5.875 0.655 ;
        RECT  5.525 0.835 5.695 1.095 ;
        RECT  5.525 2.065 5.695 3.005 ;
        RECT  5.365 0.835 5.525 3.160 ;
        RECT  4.215 3.000 5.365 3.160 ;
        RECT  5.085 0.495 5.185 1.095 ;
        RECT  5.085 2.165 5.185 2.765 ;
        RECT  4.925 0.495 5.085 2.765 ;
        RECT  4.515 0.475 4.675 2.815 ;
        RECT  4.415 0.475 4.515 0.915 ;
        RECT  4.415 2.555 4.515 2.815 ;
        RECT  3.565 0.755 4.415 0.915 ;
        RECT  4.175 1.095 4.275 1.255 ;
        RECT  4.175 2.045 4.275 2.305 ;
        RECT  4.055 2.775 4.215 3.160 ;
        RECT  4.015 1.095 4.175 2.595 ;
        RECT  2.545 2.775 4.055 2.935 ;
        RECT  2.885 2.435 4.015 2.595 ;
        RECT  3.405 0.535 3.565 1.690 ;
        RECT  2.015 0.535 3.405 0.695 ;
        RECT  3.225 2.095 3.325 2.255 ;
        RECT  3.065 0.985 3.225 2.255 ;
        RECT  2.725 1.675 2.885 2.595 ;
        RECT  2.545 0.965 2.740 1.225 ;
        RECT  2.385 0.965 2.545 2.935 ;
        RECT  1.755 0.535 2.015 1.370 ;
        RECT  1.705 2.005 1.865 2.295 ;
        RECT  1.695 1.210 1.755 1.370 ;
        RECT  1.695 2.005 1.705 2.165 ;
        RECT  1.535 1.210 1.695 2.165 ;
    END
END AHCSHCONX2

MACRO AHCSHCINX4
    CLASS CORE ;
    FOREIGN AHCSHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.585 0.695 8.615 2.810 ;
        RECT  8.415 0.695 8.585 2.920 ;
        RECT  8.325 0.695 8.415 1.295 ;
        RECT  8.325 1.980 8.415 2.920 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 2.405 7.805 2.810 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 0.485 1.915 1.085 ;
        RECT  0.895 0.925 1.655 1.085 ;
        RECT  0.945 2.275 1.205 3.215 ;
        RECT  0.335 2.275 0.945 2.435 ;
        RECT  0.580 0.485 0.895 1.085 ;
        RECT  0.270 0.925 0.580 1.085 ;
        RECT  0.270 1.700 0.335 2.435 ;
        RECT  0.110 0.925 0.270 2.435 ;
        END
        ANTENNADIFFAREA     0.9880 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.065 1.405 3.225 2.775 ;
        RECT  2.815 1.405 3.065 1.770 ;
        RECT  1.545 2.615 3.065 2.775 ;
        RECT  1.385 1.625 1.545 2.775 ;
        RECT  1.045 1.625 1.385 1.990 ;
        RECT  0.930 1.625 1.045 1.785 ;
        END
        ANTENNAGATEAREA     0.8489 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.275 1.605 2.635 1.990 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.035 -0.250 8.740 0.250 ;
        RECT  7.775 -0.250 8.035 0.405 ;
        RECT  5.025 -0.250 7.775 0.250 ;
        RECT  4.765 -0.250 5.025 0.575 ;
        RECT  2.425 -0.250 4.765 0.250 ;
        RECT  2.165 -0.250 2.425 0.740 ;
        RECT  1.405 -0.250 2.165 0.250 ;
        RECT  1.145 -0.250 1.405 0.735 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 0.735 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.035 3.440 8.740 3.940 ;
        RECT  7.775 3.285 8.035 3.940 ;
        RECT  5.155 3.440 7.775 3.940 ;
        RECT  4.895 3.115 5.155 3.940 ;
        RECT  2.395 3.440 4.895 3.940 ;
        RECT  1.795 2.955 2.395 3.940 ;
        RECT  0.385 3.440 1.795 3.940 ;
        RECT  0.125 2.615 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.075 1.535 8.235 1.795 ;
        RECT  7.945 1.535 8.075 1.695 ;
        RECT  7.785 0.675 7.945 1.695 ;
        RECT  7.435 0.675 7.785 0.835 ;
        RECT  7.555 1.035 7.605 1.295 ;
        RECT  7.555 1.955 7.605 2.215 ;
        RECT  7.345 1.035 7.555 2.215 ;
        RECT  7.275 0.495 7.435 0.835 ;
        RECT  7.125 1.525 7.345 1.785 ;
        RECT  6.585 0.495 7.275 0.655 ;
        RECT  6.945 0.835 7.095 1.095 ;
        RECT  6.945 2.045 7.095 2.985 ;
        RECT  6.835 0.835 6.945 2.985 ;
        RECT  6.785 0.835 6.835 2.205 ;
        RECT  5.495 2.825 6.835 2.985 ;
        RECT  6.485 0.495 6.585 1.095 ;
        RECT  6.485 2.045 6.585 2.645 ;
        RECT  6.325 0.495 6.485 2.645 ;
        RECT  5.975 0.755 6.075 1.015 ;
        RECT  5.975 2.045 6.075 2.645 ;
        RECT  5.815 0.755 5.975 2.645 ;
        RECT  4.585 0.755 5.815 0.915 ;
        RECT  5.120 1.095 5.565 1.255 ;
        RECT  5.120 2.035 5.565 2.295 ;
        RECT  5.335 2.775 5.495 2.985 ;
        RECT  4.065 2.775 5.335 2.935 ;
        RECT  4.960 1.095 5.120 2.595 ;
        RECT  3.905 2.435 4.960 2.595 ;
        RECT  4.585 1.415 4.775 1.675 ;
        RECT  4.245 2.095 4.605 2.255 ;
        RECT  4.425 0.485 4.585 1.675 ;
        RECT  2.935 0.485 4.425 0.645 ;
        RECT  4.085 1.040 4.245 2.255 ;
        RECT  4.005 1.040 4.085 1.200 ;
        RECT  3.565 2.775 4.065 3.035 ;
        RECT  3.745 0.940 4.005 1.200 ;
        RECT  3.745 1.575 3.905 2.595 ;
        RECT  3.405 0.940 3.565 3.035 ;
        RECT  3.185 0.940 3.405 1.200 ;
        RECT  2.675 0.485 2.935 1.085 ;
        RECT  2.725 2.170 2.885 2.430 ;
        RECT  2.035 2.170 2.725 2.330 ;
        RECT  2.470 0.925 2.675 1.085 ;
        RECT  2.310 0.925 2.470 1.425 ;
        RECT  2.085 1.265 2.310 1.425 ;
        RECT  2.035 1.265 2.085 1.525 ;
        RECT  1.875 1.265 2.035 2.330 ;
        RECT  1.825 1.265 1.875 1.525 ;
        RECT  0.450 1.265 1.825 1.425 ;
    END
END AHCSHCINX4

MACRO AHCSHCINX2
    CLASS CORE ;
    FOREIGN AHCSHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.085 0.695 7.245 3.055 ;
        RECT  6.955 0.695 7.085 1.295 ;
        RECT  7.025 2.110 7.085 3.055 ;
        RECT  6.955 2.115 7.025 3.055 ;
        END
        ANTENNADIFFAREA     0.7276 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.955 2.500 6.315 2.940 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 0.650 0.895 0.910 ;
        RECT  0.565 0.650 0.725 1.075 ;
        RECT  0.335 0.915 0.565 1.075 ;
        RECT  0.335 1.955 0.385 2.895 ;
        RECT  0.125 0.915 0.335 2.895 ;
        END
        ANTENNADIFFAREA     0.6890 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.690 2.465 1.975 2.725 ;
        RECT  0.795 2.465 1.690 2.625 ;
        RECT  0.745 1.700 0.795 2.625 ;
        RECT  0.565 1.255 0.745 2.625 ;
        RECT  0.515 1.255 0.565 1.570 ;
        END
        ANTENNAGATEAREA     0.5954 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 1.585 1.635 1.845 ;
        RECT  1.255 1.685 1.475 1.845 ;
        RECT  1.070 1.685 1.255 1.990 ;
        RECT  1.045 1.700 1.070 1.990 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.665 -0.250 7.360 0.250 ;
        RECT  6.405 -0.250 6.665 0.405 ;
        RECT  3.585 -0.250 6.405 0.250 ;
        RECT  3.325 -0.250 3.585 0.575 ;
        RECT  1.405 -0.250 3.325 0.250 ;
        RECT  1.145 -0.250 1.405 0.905 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 0.735 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.705 3.440 7.360 3.940 ;
        RECT  6.495 2.115 6.705 3.940 ;
        RECT  3.905 3.440 6.495 3.940 ;
        RECT  3.645 3.115 3.905 3.940 ;
        RECT  1.205 3.440 3.645 3.940 ;
        RECT  0.945 2.805 1.205 3.940 ;
        RECT  0.000 3.440 0.945 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.645 1.500 6.905 1.760 ;
        RECT  6.605 1.500 6.645 1.660 ;
        RECT  6.445 0.675 6.605 1.660 ;
        RECT  6.055 0.675 6.445 0.835 ;
        RECT  6.015 1.035 6.225 1.435 ;
        RECT  6.015 1.955 6.115 2.215 ;
        RECT  5.895 0.495 6.055 0.835 ;
        RECT  5.965 1.035 6.015 2.215 ;
        RECT  5.855 1.275 5.965 2.215 ;
        RECT  5.205 0.495 5.895 0.655 ;
        RECT  5.765 1.525 5.855 1.785 ;
        RECT  5.585 0.835 5.715 1.095 ;
        RECT  5.585 2.465 5.715 2.725 ;
        RECT  5.425 0.835 5.585 3.140 ;
        RECT  4.245 2.980 5.425 3.140 ;
        RECT  5.165 0.495 5.205 1.095 ;
        RECT  5.165 2.110 5.205 2.710 ;
        RECT  5.005 0.495 5.165 2.710 ;
        RECT  4.945 0.495 5.005 1.095 ;
        RECT  4.945 2.110 5.005 2.710 ;
        RECT  4.645 0.755 4.695 1.020 ;
        RECT  4.645 2.540 4.695 2.800 ;
        RECT  4.485 0.755 4.645 2.800 ;
        RECT  4.435 0.755 4.485 1.020 ;
        RECT  4.435 2.540 4.485 2.800 ;
        RECT  3.475 0.755 4.435 0.915 ;
        RECT  4.195 2.030 4.295 2.290 ;
        RECT  4.085 2.775 4.245 3.140 ;
        RECT  4.035 1.095 4.195 2.595 ;
        RECT  2.770 2.775 4.085 2.935 ;
        RECT  3.920 1.095 4.035 1.255 ;
        RECT  2.655 2.435 4.035 2.595 ;
        RECT  3.475 1.425 3.525 1.685 ;
        RECT  3.265 0.755 3.475 1.685 ;
        RECT  2.995 2.095 3.355 2.255 ;
        RECT  2.965 0.755 3.265 0.915 ;
        RECT  2.835 1.095 2.995 2.255 ;
        RECT  2.805 0.545 2.965 0.915 ;
        RECT  2.735 1.095 2.835 1.255 ;
        RECT  1.975 0.545 2.805 0.705 ;
        RECT  2.510 2.775 2.770 3.035 ;
        RECT  2.495 1.585 2.655 2.595 ;
        RECT  2.315 2.775 2.510 2.935 ;
        RECT  2.315 0.905 2.485 1.165 ;
        RECT  2.225 0.905 2.315 2.935 ;
        RECT  2.155 1.005 2.225 2.935 ;
        RECT  1.815 0.545 1.975 2.185 ;
        RECT  1.715 0.545 1.815 1.365 ;
        RECT  1.715 2.025 1.815 2.185 ;
        RECT  1.235 1.205 1.715 1.365 ;
        RECT  1.455 2.025 1.715 2.285 ;
        RECT  0.945 1.205 1.235 1.465 ;
    END
END AHCSHCINX2

MACRO ACCSIHCONX4
    CLASS CORE ;
    FOREIGN ACCSIHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.215 0.855 4.475 2.435 ;
        RECT  2.505 0.855 4.215 1.115 ;
        RECT  3.300 2.175 4.215 2.435 ;
        RECT  3.040 2.175 3.300 3.135 ;
        END
        ANTENNADIFFAREA     1.0660 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 2.290 1.915 2.890 ;
        RECT  0.895 2.290 1.655 2.450 ;
        RECT  0.945 0.515 1.205 1.115 ;
        RECT  0.725 0.880 0.945 1.115 ;
        RECT  0.585 2.290 0.895 2.890 ;
        RECT  0.565 0.880 0.725 1.495 ;
        RECT  0.335 2.290 0.585 2.450 ;
        RECT  0.335 1.335 0.565 1.495 ;
        RECT  0.130 1.335 0.335 2.450 ;
        RECT  0.125 1.335 0.130 2.400 ;
        END
        ANTENNADIFFAREA     1.0564 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.725 1.295 3.985 1.665 ;
        RECT  2.595 1.295 3.725 1.455 ;
        RECT  2.265 1.295 2.595 1.625 ;
        RECT  2.150 1.295 2.265 1.580 ;
        RECT  1.715 1.295 2.150 1.455 ;
        RECT  1.505 1.290 1.715 1.580 ;
        RECT  1.375 1.295 1.505 1.580 ;
        RECT  1.165 1.295 1.375 1.675 ;
        RECT  1.115 1.415 1.165 1.675 ;
        END
        ANTENNAGATEAREA     0.9802 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 1.635 3.475 1.795 ;
        RECT  2.775 1.635 2.935 1.995 ;
        RECT  2.635 1.835 2.775 1.995 ;
        RECT  2.425 1.835 2.635 2.400 ;
        RECT  2.085 1.835 2.425 2.015 ;
        RECT  1.985 1.775 2.085 2.015 ;
        RECT  1.825 1.775 1.985 2.020 ;
        RECT  0.675 1.860 1.825 2.020 ;
        RECT  0.515 1.725 0.675 2.020 ;
        END
        ANTENNAGATEAREA     0.9802 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 -0.250 4.600 0.250 ;
        RECT  4.125 -0.250 4.385 0.405 ;
        RECT  3.305 -0.250 4.125 0.250 ;
        RECT  3.045 -0.250 3.305 0.405 ;
        RECT  2.085 -0.250 3.045 0.250 ;
        RECT  1.825 -0.250 2.085 1.075 ;
        RECT  0.385 -0.250 1.825 0.250 ;
        RECT  0.125 -0.250 0.385 1.075 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.155 3.440 4.600 3.940 ;
        RECT  3.895 2.615 4.155 3.940 ;
        RECT  2.455 3.440 3.895 3.940 ;
        RECT  2.195 2.590 2.455 3.940 ;
        RECT  1.405 3.440 2.195 3.940 ;
        RECT  1.145 2.755 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.755 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END ACCSIHCONX4

MACRO ACCSIHCONX2
    CLASS CORE ;
    FOREIGN ACCSIHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.575 2.255 2.895 ;
        RECT  1.815 1.575 1.965 1.835 ;
        RECT  1.555 0.750 1.815 1.835 ;
        RECT  1.485 0.750 1.555 1.010 ;
        END
        ANTENNADIFFAREA     0.6890 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.110 1.715 2.400 ;
        RECT  1.375 2.110 1.505 2.330 ;
        RECT  1.215 1.245 1.375 2.330 ;
        RECT  0.745 1.245 1.215 1.405 ;
        RECT  0.895 2.170 1.215 2.330 ;
        RECT  0.635 2.170 0.895 2.770 ;
        RECT  0.585 1.035 0.745 1.405 ;
        RECT  0.385 1.035 0.585 1.195 ;
        RECT  0.125 0.595 0.385 1.195 ;
        END
        ANTENNADIFFAREA     0.6572 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.475 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.4901 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.745 1.585 1.035 1.990 ;
        RECT  0.585 1.700 0.745 1.990 ;
        END
        ANTENNAGATEAREA     0.4901 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.255 -0.250 2.760 0.250 ;
        RECT  1.995 -0.250 2.255 1.285 ;
        RECT  1.205 -0.250 1.995 0.250 ;
        RECT  0.945 -0.250 1.205 1.060 ;
        RECT  0.000 -0.250 0.945 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 3.440 2.760 3.940 ;
        RECT  1.175 2.615 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END ACCSIHCONX2

MACRO ACCSHCONX4
    CLASS CORE ;
    FOREIGN ACCSHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.040 0.810 9.300 1.240 ;
        RECT  8.190 0.810 9.040 0.970 ;
        RECT  8.805 2.080 8.995 2.240 ;
        RECT  8.645 2.025 8.805 2.240 ;
        RECT  8.155 2.025 8.645 2.185 ;
        RECT  8.155 0.810 8.190 1.295 ;
        RECT  8.030 0.810 8.155 2.185 ;
        RECT  8.005 1.035 8.030 2.185 ;
        RECT  7.930 1.035 8.005 2.305 ;
        RECT  7.875 2.025 7.930 2.305 ;
        RECT  7.715 2.025 7.875 2.540 ;
        RECT  6.995 2.380 7.715 2.540 ;
        RECT  6.995 0.695 7.170 1.295 ;
        RECT  6.910 0.695 6.995 2.540 ;
        RECT  6.835 1.135 6.910 2.540 ;
        RECT  6.665 2.105 6.835 2.400 ;
        END
        ANTENNADIFFAREA     1.8301 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.780 2.275 12.040 3.215 ;
        RECT  10.935 3.050 11.780 3.210 ;
        RECT  10.915 1.150 11.340 1.310 ;
        RECT  10.915 2.405 10.935 3.210 ;
        RECT  10.705 1.150 10.915 3.210 ;
        RECT  10.320 1.150 10.705 1.360 ;
        RECT  10.675 2.405 10.705 3.210 ;
        RECT  10.390 3.050 10.675 3.210 ;
        RECT  10.230 3.050 10.390 3.260 ;
        RECT  10.060 0.810 10.320 1.360 ;
        RECT  9.625 3.100 10.230 3.260 ;
        END
        ANTENNADIFFAREA     1.8130 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.135 1.470 14.340 1.730 ;
        RECT  13.925 1.470 14.135 1.990 ;
        RECT  13.740 1.470 13.925 1.730 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.205 1.290 13.215 1.580 ;
        RECT  13.005 1.290 13.205 1.675 ;
        RECT  12.265 1.415 13.005 1.675 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 1.515 5.045 1.775 ;
        RECT  4.725 1.515 4.935 1.990 ;
        RECT  4.445 1.515 4.725 1.775 ;
        END
        ANTENNAGATEAREA     0.8268 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.515 0.455 1.915 ;
        RECT  0.125 1.515 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.595 -0.250 14.720 0.250 ;
        RECT  14.335 -0.250 14.595 1.195 ;
        RECT  13.535 -0.250 14.335 0.250 ;
        RECT  12.595 -0.250 13.535 0.405 ;
        RECT  6.605 -0.250 12.595 0.250 ;
        RECT  6.005 -0.250 6.605 1.135 ;
        RECT  4.815 -0.250 6.005 0.250 ;
        RECT  4.555 -0.250 4.815 1.195 ;
        RECT  1.835 -0.250 4.555 0.250 ;
        RECT  1.575 -0.250 1.835 0.405 ;
        RECT  0.385 -0.250 1.575 0.250 ;
        RECT  0.125 -0.250 0.385 1.195 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.595 3.440 14.720 3.940 ;
        RECT  14.335 2.105 14.595 3.940 ;
        RECT  13.575 3.440 14.335 3.940 ;
        RECT  13.315 2.535 13.575 3.940 ;
        RECT  12.555 3.440 13.315 3.940 ;
        RECT  12.295 2.255 12.555 3.940 ;
        RECT  5.875 3.440 12.295 3.940 ;
        RECT  5.615 3.285 5.875 3.940 ;
        RECT  4.845 3.440 5.615 3.940 ;
        RECT  4.585 3.285 4.845 3.940 ;
        RECT  1.835 3.440 4.585 3.940 ;
        RECT  1.575 3.285 1.835 3.940 ;
        RECT  0.385 3.440 1.575 3.940 ;
        RECT  0.125 2.250 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.825 0.585 14.085 1.195 ;
        RECT  13.825 2.170 14.085 3.110 ;
        RECT  12.285 0.585 13.825 0.745 ;
        RECT  13.555 1.035 13.825 1.195 ;
        RECT  13.555 2.170 13.825 2.330 ;
        RECT  13.395 1.035 13.555 2.330 ;
        RECT  12.805 1.910 13.065 3.080 ;
        RECT  11.885 0.930 12.990 1.090 ;
        RECT  11.885 1.910 12.805 2.070 ;
        RECT  12.125 0.470 12.285 0.745 ;
        RECT  7.680 0.470 12.125 0.630 ;
        RECT  11.880 0.930 11.885 2.070 ;
        RECT  11.725 0.810 11.880 2.070 ;
        RECT  11.620 0.810 11.725 1.140 ;
        RECT  11.530 1.910 11.725 2.070 ;
        RECT  10.570 0.810 11.620 0.970 ;
        RECT  11.270 1.910 11.530 2.625 ;
        RECT  9.810 2.490 10.425 2.750 ;
        RECT  9.650 0.810 9.810 2.920 ;
        RECT  9.550 0.810 9.650 1.360 ;
        RECT  9.445 2.760 9.650 2.920 ;
        RECT  9.285 2.760 9.445 3.220 ;
        RECT  9.175 1.490 9.335 2.580 ;
        RECT  6.220 3.060 9.285 3.220 ;
        RECT  8.735 1.490 9.175 1.650 ;
        RECT  8.485 2.420 9.175 2.580 ;
        RECT  8.735 1.150 8.790 1.310 ;
        RECT  8.575 1.150 8.735 1.650 ;
        RECT  8.530 1.150 8.575 1.310 ;
        RECT  8.385 2.370 8.485 2.630 ;
        RECT  8.225 2.370 8.385 2.880 ;
        RECT  6.600 2.720 8.225 2.880 ;
        RECT  7.580 0.470 7.680 1.195 ;
        RECT  7.465 0.470 7.580 1.800 ;
        RECT  7.420 0.470 7.465 2.200 ;
        RECT  7.305 1.640 7.420 2.200 ;
        RECT  7.175 2.040 7.305 2.200 ;
        RECT  6.365 1.315 6.615 1.475 ;
        RECT  6.440 2.600 6.600 2.880 ;
        RECT  6.005 2.600 6.440 2.760 ;
        RECT  6.205 1.315 6.365 2.215 ;
        RECT  6.060 2.945 6.220 3.220 ;
        RECT  5.725 1.315 6.205 1.475 ;
        RECT  4.355 2.945 6.060 3.105 ;
        RECT  5.845 2.055 6.005 2.760 ;
        RECT  5.385 2.055 5.845 2.215 ;
        RECT  5.565 0.495 5.725 1.475 ;
        RECT  3.905 2.395 5.645 2.555 ;
        RECT  5.465 0.495 5.565 0.755 ;
        RECT  5.225 1.035 5.385 2.215 ;
        RECT  5.065 1.035 5.225 1.295 ;
        RECT  5.125 1.955 5.225 2.215 ;
        RECT  4.195 2.945 4.355 3.190 ;
        RECT  4.255 0.495 4.305 0.755 ;
        RECT  4.255 1.955 4.305 2.215 ;
        RECT  4.095 0.495 4.255 2.215 ;
        RECT  2.265 3.030 4.195 3.190 ;
        RECT  4.045 0.495 4.095 0.755 ;
        RECT  4.045 1.955 4.095 2.215 ;
        RECT  3.425 0.585 4.045 0.745 ;
        RECT  3.805 1.035 3.905 1.295 ;
        RECT  3.805 2.395 3.905 2.840 ;
        RECT  3.645 1.035 3.805 2.840 ;
        RECT  2.885 2.680 3.645 2.840 ;
        RECT  3.245 0.955 3.395 1.215 ;
        RECT  3.245 2.340 3.395 2.500 ;
        RECT  3.085 0.585 3.245 2.500 ;
        RECT  1.300 0.585 3.085 0.745 ;
        RECT  2.725 0.925 2.885 2.840 ;
        RECT  2.625 0.925 2.725 1.185 ;
        RECT  2.625 2.465 2.725 2.840 ;
        RECT  2.215 0.925 2.375 2.640 ;
        RECT  2.105 2.945 2.265 3.190 ;
        RECT  2.115 0.925 2.215 1.185 ;
        RECT  2.115 2.040 2.215 2.640 ;
        RECT  0.795 2.945 2.105 3.105 ;
        RECT  1.300 1.585 2.035 1.845 ;
        RECT  1.235 0.585 1.300 1.845 ;
        RECT  1.235 2.480 1.295 2.740 ;
        RECT  1.140 0.585 1.235 2.740 ;
        RECT  1.075 1.035 1.140 2.740 ;
        RECT  1.035 1.035 1.075 1.295 ;
        RECT  1.035 2.480 1.075 2.740 ;
        RECT  0.795 0.495 0.895 0.755 ;
        RECT  0.795 1.955 0.895 2.215 ;
        RECT  0.635 0.495 0.795 3.105 ;
    END
END ACCSHCONX4

MACRO ACCSHCONX2
    CLASS CORE ;
    FOREIGN ACCSHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.385 0.810 8.645 1.240 ;
        RECT  8.345 2.080 8.455 2.240 ;
        RECT  7.565 0.810 8.385 0.970 ;
        RECT  8.185 1.830 8.345 2.240 ;
        RECT  7.695 1.830 8.185 1.990 ;
        RECT  7.465 1.700 7.695 1.990 ;
        RECT  7.465 0.810 7.565 1.295 ;
        RECT  7.435 0.810 7.465 2.185 ;
        RECT  7.405 0.810 7.435 2.410 ;
        RECT  7.305 1.035 7.405 2.410 ;
        RECT  7.175 2.025 7.305 2.410 ;
        END
        ANTENNADIFFAREA     1.0759 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.055 0.810 10.185 1.860 ;
        RECT  10.055 2.405 10.155 3.005 ;
        RECT  10.025 0.810 10.055 3.210 ;
        RECT  9.155 0.810 10.025 0.970 ;
        RECT  9.895 1.700 10.025 3.210 ;
        RECT  9.785 1.700 9.895 1.990 ;
        RECT  9.785 3.050 9.895 3.210 ;
        RECT  9.450 3.050 9.785 3.260 ;
        RECT  8.845 3.100 9.450 3.260 ;
        RECT  8.895 0.810 9.155 1.240 ;
        END
        ANTENNADIFFAREA     1.1482 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.520 1.515 11.835 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.705 1.290 11.000 1.800 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 1.515 5.045 1.775 ;
        RECT  4.725 1.515 4.935 1.990 ;
        RECT  4.445 1.515 4.725 1.775 ;
        END
        ANTENNAGATEAREA     0.8268 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.515 0.455 1.915 ;
        RECT  0.125 1.515 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.295 -0.250 11.960 0.250 ;
        RECT  11.035 -0.250 11.295 0.405 ;
        RECT  6.375 -0.250 11.035 0.250 ;
        RECT  6.115 -0.250 6.375 1.135 ;
        RECT  6.055 -0.250 6.115 0.405 ;
        RECT  4.815 -0.250 6.055 0.250 ;
        RECT  4.555 -0.250 4.815 1.195 ;
        RECT  1.835 -0.250 4.555 0.250 ;
        RECT  1.575 -0.250 1.835 0.405 ;
        RECT  0.385 -0.250 1.575 0.250 ;
        RECT  0.125 -0.250 0.385 1.195 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.255 3.440 11.960 3.940 ;
        RECT  10.995 2.535 11.255 3.940 ;
        RECT  5.875 3.440 10.995 3.940 ;
        RECT  5.615 3.285 5.875 3.940 ;
        RECT  4.845 3.440 5.615 3.940 ;
        RECT  4.585 3.285 4.845 3.940 ;
        RECT  1.835 3.440 4.585 3.940 ;
        RECT  1.575 3.285 1.835 3.940 ;
        RECT  0.385 3.440 1.575 3.940 ;
        RECT  0.125 2.250 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.575 0.585 11.835 1.195 ;
        RECT  11.575 2.170 11.835 3.110 ;
        RECT  10.720 0.585 11.575 0.745 ;
        RECT  11.340 1.035 11.575 1.195 ;
        RECT  11.340 2.170 11.575 2.330 ;
        RECT  11.180 1.035 11.340 2.330 ;
        RECT  10.525 0.935 10.755 1.095 ;
        RECT  10.560 0.470 10.720 0.745 ;
        RECT  10.525 2.140 10.665 3.080 ;
        RECT  7.055 0.470 10.560 0.630 ;
        RECT  10.405 0.935 10.525 3.080 ;
        RECT  10.365 0.935 10.405 2.300 ;
        RECT  9.595 1.150 9.695 1.310 ;
        RECT  9.595 2.490 9.645 2.750 ;
        RECT  9.435 1.150 9.595 2.750 ;
        RECT  9.385 2.490 9.435 2.750 ;
        RECT  9.135 2.590 9.385 2.750 ;
        RECT  8.975 2.590 9.135 2.920 ;
        RECT  8.300 2.760 8.975 2.920 ;
        RECT  8.635 1.490 8.795 2.580 ;
        RECT  8.195 1.490 8.635 1.650 ;
        RECT  7.945 2.420 8.635 2.580 ;
        RECT  8.140 2.760 8.300 3.110 ;
        RECT  8.035 1.150 8.195 1.650 ;
        RECT  6.215 2.950 8.140 3.110 ;
        RECT  7.845 1.150 8.035 1.310 ;
        RECT  7.685 2.370 7.945 2.760 ;
        RECT  5.995 2.600 7.685 2.760 ;
        RECT  6.955 0.470 7.055 1.295 ;
        RECT  6.895 0.470 6.955 2.305 ;
        RECT  6.795 1.035 6.895 2.305 ;
        RECT  6.665 2.045 6.795 2.305 ;
        RECT  6.365 1.315 6.615 1.475 ;
        RECT  6.205 1.315 6.365 2.215 ;
        RECT  6.055 2.945 6.215 3.110 ;
        RECT  5.775 1.315 6.205 1.505 ;
        RECT  4.260 2.945 6.055 3.105 ;
        RECT  5.835 2.055 5.995 2.760 ;
        RECT  5.385 2.055 5.835 2.215 ;
        RECT  5.615 0.495 5.775 1.505 ;
        RECT  3.905 2.395 5.645 2.555 ;
        RECT  5.515 0.495 5.615 0.755 ;
        RECT  5.225 1.035 5.385 2.215 ;
        RECT  5.065 1.035 5.225 1.295 ;
        RECT  5.125 1.955 5.225 2.215 ;
        RECT  4.255 0.495 4.305 0.755 ;
        RECT  4.255 1.955 4.305 2.215 ;
        RECT  4.100 2.945 4.260 3.190 ;
        RECT  4.095 0.495 4.255 2.215 ;
        RECT  2.260 3.030 4.100 3.190 ;
        RECT  4.045 0.495 4.095 0.755 ;
        RECT  4.045 1.955 4.095 2.215 ;
        RECT  3.425 0.585 4.045 0.745 ;
        RECT  3.805 1.035 3.905 1.295 ;
        RECT  3.805 2.395 3.905 2.840 ;
        RECT  3.645 1.035 3.805 2.840 ;
        RECT  2.885 2.680 3.645 2.840 ;
        RECT  3.245 0.955 3.395 1.215 ;
        RECT  3.245 2.340 3.395 2.500 ;
        RECT  3.085 0.585 3.245 2.500 ;
        RECT  1.300 0.585 3.085 0.745 ;
        RECT  2.725 0.925 2.885 2.840 ;
        RECT  2.625 0.925 2.725 1.185 ;
        RECT  2.625 2.465 2.725 2.725 ;
        RECT  2.215 0.925 2.375 2.640 ;
        RECT  2.100 2.945 2.260 3.190 ;
        RECT  2.115 0.925 2.215 1.185 ;
        RECT  2.115 2.040 2.215 2.640 ;
        RECT  0.795 2.945 2.100 3.105 ;
        RECT  1.300 1.585 2.035 1.845 ;
        RECT  1.235 0.585 1.300 1.845 ;
        RECT  1.235 2.480 1.295 2.740 ;
        RECT  1.140 0.585 1.235 2.740 ;
        RECT  1.075 1.035 1.140 2.740 ;
        RECT  1.035 1.035 1.075 1.295 ;
        RECT  1.035 2.480 1.075 2.740 ;
        RECT  0.795 0.495 0.895 0.755 ;
        RECT  0.795 1.955 0.895 2.215 ;
        RECT  0.635 0.495 0.795 3.105 ;
    END
END ACCSHCONX2

MACRO ACCSHCINX4
    CLASS CORE ;
    FOREIGN ACCSHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.615 1.015 11.775 1.860 ;
        RECT  10.915 1.700 11.615 1.860 ;
        RECT  10.915 2.280 11.125 2.540 ;
        RECT  10.705 1.700 10.915 2.540 ;
        RECT  10.545 0.565 10.805 1.165 ;
        RECT  9.285 2.380 10.705 2.540 ;
        RECT  10.185 1.005 10.545 1.165 ;
        RECT  10.025 1.005 10.185 1.830 ;
        RECT  9.285 1.670 10.025 1.830 ;
        RECT  9.125 1.670 9.285 2.540 ;
        RECT  8.925 1.920 9.125 2.080 ;
        END
        ANTENNADIFFAREA     2.0685 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.490 1.265 14.465 1.425 ;
        RECT  14.145 2.405 14.405 3.015 ;
        RECT  13.385 2.855 14.145 3.015 ;
        RECT  13.415 1.265 13.490 1.580 ;
        RECT  13.385 1.015 13.415 1.580 ;
        RECT  13.225 1.015 13.385 3.015 ;
        RECT  13.155 1.015 13.225 1.275 ;
        RECT  13.005 2.110 13.225 3.015 ;
        RECT  12.365 2.855 13.005 3.015 ;
        RECT  12.105 2.745 12.365 3.015 ;
        END
        ANTENNADIFFAREA     1.5015 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.145 1.635 16.505 1.990 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.195 1.585 15.550 1.990 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.540 1.245 7.335 1.405 ;
        RECT  6.490 0.810 6.540 1.405 ;
        RECT  6.330 0.810 6.490 2.055 ;
        RECT  6.280 0.810 6.330 1.170 ;
        RECT  6.290 1.700 6.330 2.055 ;
        RECT  6.150 1.895 6.290 2.055 ;
        RECT  6.105 0.880 6.280 1.170 ;
        RECT  5.990 1.895 6.150 2.155 ;
        END
        ANTENNAGATEAREA     0.8268 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.430 0.440 1.985 ;
        RECT  0.125 1.430 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.355 -0.250 17.480 0.250 ;
        RECT  17.095 -0.250 17.355 1.190 ;
        RECT  16.335 -0.250 17.095 0.250 ;
        RECT  16.075 -0.250 16.335 1.095 ;
        RECT  15.015 -0.250 16.075 0.250 ;
        RECT  14.755 -0.250 15.015 0.405 ;
        RECT  9.990 -0.250 14.755 0.250 ;
        RECT  9.730 -0.250 9.990 0.405 ;
        RECT  8.670 -0.250 9.730 0.250 ;
        RECT  8.410 -0.250 8.670 0.405 ;
        RECT  7.520 -0.250 8.410 0.250 ;
        RECT  7.260 -0.250 7.520 0.405 ;
        RECT  1.010 -0.250 7.260 0.250 ;
        RECT  0.750 -0.250 1.010 0.405 ;
        RECT  0.000 -0.250 0.750 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.355 3.440 17.480 3.940 ;
        RECT  17.095 2.255 17.355 3.940 ;
        RECT  16.335 3.440 17.095 3.940 ;
        RECT  16.075 2.255 16.335 3.940 ;
        RECT  15.315 3.440 16.075 3.940 ;
        RECT  15.055 2.935 15.315 3.940 ;
        RECT  7.780 3.440 15.055 3.940 ;
        RECT  7.520 3.285 7.780 3.940 ;
        RECT  1.835 3.440 7.520 3.940 ;
        RECT  1.575 3.285 1.835 3.940 ;
        RECT  0.385 3.440 1.575 3.940 ;
        RECT  0.125 2.255 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.685 0.695 16.845 3.195 ;
        RECT  16.585 0.695 16.685 1.450 ;
        RECT  16.585 2.255 16.685 3.195 ;
        RECT  15.895 1.290 16.585 1.450 ;
        RECT  15.735 0.585 15.895 1.450 ;
        RECT  15.565 2.255 15.825 3.195 ;
        RECT  14.340 0.585 15.735 0.745 ;
        RECT  14.920 2.255 15.565 2.470 ;
        RECT  15.295 0.925 15.555 1.185 ;
        RECT  14.920 0.925 15.295 1.085 ;
        RECT  14.915 0.925 14.920 2.470 ;
        RECT  14.760 0.925 14.915 2.595 ;
        RECT  13.925 0.925 14.760 1.085 ;
        RECT  14.655 2.065 14.760 2.595 ;
        RECT  13.895 2.065 14.655 2.225 ;
        RECT  14.180 0.470 14.340 0.745 ;
        RECT  11.315 0.470 14.180 0.630 ;
        RECT  13.665 0.825 13.925 1.085 ;
        RECT  13.735 2.065 13.895 2.510 ;
        RECT  13.635 2.250 13.735 2.510 ;
        RECT  12.825 0.810 12.975 1.920 ;
        RECT  12.815 0.810 12.825 2.665 ;
        RECT  12.115 0.810 12.815 0.970 ;
        RECT  12.665 1.760 12.815 2.665 ;
        RECT  12.295 1.270 12.455 2.555 ;
        RECT  11.805 2.395 12.295 2.555 ;
        RECT  11.955 0.810 12.115 2.205 ;
        RECT  11.465 2.045 11.955 2.205 ;
        RECT  11.645 2.395 11.805 3.220 ;
        RECT  8.515 3.060 11.645 3.220 ;
        RECT  11.305 2.045 11.465 2.880 ;
        RECT  11.215 0.470 11.315 1.175 ;
        RECT  8.945 2.720 11.305 2.880 ;
        RECT  11.055 0.470 11.215 1.505 ;
        RECT  10.525 1.345 11.055 1.505 ;
        RECT  10.365 1.345 10.525 2.170 ;
        RECT  7.080 0.585 10.365 0.745 ;
        RECT  9.465 2.010 10.365 2.170 ;
        RECT  8.490 0.945 9.415 1.105 ;
        RECT  8.785 2.265 8.945 2.880 ;
        RECT  6.995 2.265 8.785 2.425 ;
        RECT  7.000 2.605 8.605 2.765 ;
        RECT  8.355 2.945 8.515 3.220 ;
        RECT  8.330 0.945 8.490 2.085 ;
        RECT  7.340 2.945 8.355 3.105 ;
        RECT  7.275 1.925 8.330 2.085 ;
        RECT  8.000 0.925 8.100 1.085 ;
        RECT  7.840 0.925 8.000 1.745 ;
        RECT  6.995 1.585 7.840 1.745 ;
        RECT  7.180 2.945 7.340 3.220 ;
        RECT  2.175 3.060 7.180 3.220 ;
        RECT  6.920 0.470 7.080 0.745 ;
        RECT  6.840 2.605 7.000 2.880 ;
        RECT  6.835 1.585 6.995 2.425 ;
        RECT  5.925 0.470 6.920 0.630 ;
        RECT  2.515 2.720 6.840 2.880 ;
        RECT  6.585 2.255 6.835 2.425 ;
        RECT  6.420 2.255 6.585 2.495 ;
        RECT  6.250 2.335 6.420 2.495 ;
        RECT  5.805 2.380 5.965 2.540 ;
        RECT  5.805 0.470 5.925 1.715 ;
        RECT  5.765 0.470 5.805 2.540 ;
        RECT  5.125 0.470 5.765 0.630 ;
        RECT  5.645 1.555 5.765 2.540 ;
        RECT  5.455 0.930 5.585 1.375 ;
        RECT  5.425 0.930 5.455 2.540 ;
        RECT  5.295 1.215 5.425 2.540 ;
        RECT  2.855 2.380 5.295 2.540 ;
        RECT  5.025 0.470 5.125 1.020 ;
        RECT  4.965 0.470 5.025 2.165 ;
        RECT  4.865 0.760 4.965 2.165 ;
        RECT  4.655 2.005 4.865 2.165 ;
        RECT  4.405 0.470 4.615 1.195 ;
        RECT  4.245 0.470 4.405 2.200 ;
        RECT  3.235 0.470 4.245 0.785 ;
        RECT  3.165 2.040 4.245 2.200 ;
        RECT  2.915 1.035 3.935 1.295 ;
        RECT  1.595 0.470 3.235 0.630 ;
        RECT  2.655 0.810 2.915 1.295 ;
        RECT  2.695 2.245 2.855 2.540 ;
        RECT  2.275 2.245 2.695 2.405 ;
        RECT  1.935 0.810 2.655 0.970 ;
        RECT  2.355 2.605 2.515 2.880 ;
        RECT  2.275 1.150 2.375 1.310 ;
        RECT  1.935 2.605 2.355 2.765 ;
        RECT  2.115 1.150 2.275 2.405 ;
        RECT  2.015 2.945 2.175 3.220 ;
        RECT  1.595 2.945 2.015 3.105 ;
        RECT  1.775 0.810 1.935 2.765 ;
        RECT  1.435 0.470 1.595 0.755 ;
        RECT  1.435 1.135 1.595 3.105 ;
        RECT  0.385 0.595 1.435 0.755 ;
        RECT  1.425 1.135 1.435 1.295 ;
        RECT  1.295 2.935 1.435 3.105 ;
        RECT  1.165 1.035 1.425 1.295 ;
        RECT  1.035 2.935 1.295 3.195 ;
        RECT  0.895 1.570 1.255 1.830 ;
        RECT  0.635 1.035 0.895 2.555 ;
        RECT  0.385 1.035 0.635 1.195 ;
        RECT  0.125 0.595 0.385 1.195 ;
    END
END ACCSHCINX4

MACRO ACCSHCINX2
    CLASS CORE ;
    FOREIGN ACCSHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.385 0.885 10.545 2.540 ;
        RECT  10.375 0.885 10.385 2.510 ;
        RECT  10.245 1.700 10.375 2.510 ;
        RECT  9.995 1.700 10.245 1.925 ;
        RECT  9.050 2.350 10.245 2.510 ;
        RECT  9.785 1.700 9.995 1.990 ;
        RECT  8.890 1.920 9.050 2.510 ;
        RECT  8.650 1.920 8.890 2.080 ;
        END
        ANTENNADIFFAREA     1.2598 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.890 2.510 13.065 3.110 ;
        RECT  12.890 0.915 13.005 1.175 ;
        RECT  12.730 0.915 12.890 3.110 ;
        RECT  12.545 1.355 12.730 1.990 ;
        RECT  12.015 2.855 12.730 3.015 ;
        RECT  11.905 1.355 12.545 1.515 ;
        RECT  11.755 2.745 12.015 3.015 ;
        RECT  11.745 1.150 11.905 1.515 ;
        END
        ANTENNADIFFAREA     1.1773 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.925 1.290 14.255 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.525 1.365 13.745 1.990 ;
        RECT  13.465 1.700 13.525 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 1.245 7.225 1.405 ;
        RECT  6.385 0.810 6.435 1.405 ;
        RECT  6.175 0.810 6.385 2.055 ;
        RECT  6.150 0.880 6.175 2.055 ;
        RECT  6.105 0.880 6.150 2.155 ;
        RECT  5.990 1.895 6.105 2.155 ;
        END
        ANTENNAGATEAREA     0.8268 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.430 0.440 1.985 ;
        RECT  0.125 1.430 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.055 -0.250 14.720 0.250 ;
        RECT  13.795 -0.250 14.055 0.405 ;
        RECT  9.445 -0.250 13.795 0.250 ;
        RECT  9.185 -0.250 9.445 0.405 ;
        RECT  8.475 -0.250 9.185 0.250 ;
        RECT  8.215 -0.250 8.475 0.405 ;
        RECT  7.325 -0.250 8.215 0.250 ;
        RECT  7.065 -0.250 7.325 0.405 ;
        RECT  1.010 -0.250 7.065 0.250 ;
        RECT  0.750 -0.250 1.010 0.405 ;
        RECT  0.000 -0.250 0.750 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.085 3.440 14.720 3.940 ;
        RECT  13.825 2.255 14.085 3.940 ;
        RECT  7.780 3.440 13.825 3.940 ;
        RECT  7.520 3.285 7.780 3.940 ;
        RECT  1.835 3.440 7.520 3.940 ;
        RECT  1.575 3.285 1.835 3.940 ;
        RECT  0.385 3.440 1.575 3.940 ;
        RECT  0.125 2.255 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.435 0.495 14.595 3.195 ;
        RECT  14.335 0.495 14.435 1.095 ;
        RECT  14.335 2.255 14.435 3.195 ;
        RECT  13.405 0.585 14.335 0.745 ;
        RECT  13.315 2.170 13.575 3.195 ;
        RECT  13.345 0.925 13.515 1.185 ;
        RECT  13.245 0.470 13.405 0.745 ;
        RECT  13.285 0.925 13.345 1.520 ;
        RECT  13.285 2.170 13.315 2.330 ;
        RECT  13.185 0.925 13.285 2.330 ;
        RECT  10.155 0.470 13.245 0.630 ;
        RECT  13.125 1.360 13.185 2.330 ;
        RECT  12.425 2.405 12.525 2.665 ;
        RECT  12.235 0.810 12.495 1.175 ;
        RECT  12.265 2.230 12.425 2.665 ;
        RECT  11.565 2.230 12.265 2.390 ;
        RECT  11.565 0.810 12.235 0.970 ;
        RECT  11.405 0.810 11.565 2.390 ;
        RECT  10.885 0.810 11.405 0.970 ;
        RECT  11.065 1.270 11.225 3.220 ;
        RECT  8.125 3.060 11.065 3.220 ;
        RECT  10.725 0.810 10.885 2.880 ;
        RECT  8.710 2.720 10.725 2.880 ;
        RECT  10.075 0.470 10.155 1.225 ;
        RECT  9.995 0.470 10.075 1.275 ;
        RECT  9.975 1.015 9.995 1.275 ;
        RECT  9.815 1.015 9.975 1.505 ;
        RECT  6.825 0.585 9.815 0.745 ;
        RECT  9.510 1.345 9.815 1.505 ;
        RECT  9.350 1.345 9.510 2.165 ;
        RECT  9.230 2.005 9.350 2.165 ;
        RECT  8.245 0.945 9.045 1.105 ;
        RECT  8.550 2.265 8.710 2.880 ;
        RECT  6.800 2.265 8.550 2.425 ;
        RECT  7.000 2.605 8.370 2.765 ;
        RECT  8.085 0.945 8.245 2.085 ;
        RECT  7.965 2.945 8.125 3.220 ;
        RECT  7.275 1.925 8.085 2.085 ;
        RECT  7.340 2.945 7.965 3.105 ;
        RECT  7.805 0.925 7.905 1.085 ;
        RECT  7.645 0.925 7.805 1.745 ;
        RECT  6.800 1.585 7.645 1.745 ;
        RECT  7.180 2.945 7.340 3.220 ;
        RECT  2.175 3.060 7.180 3.220 ;
        RECT  6.840 2.605 7.000 2.880 ;
        RECT  2.515 2.720 6.840 2.880 ;
        RECT  6.665 0.470 6.825 0.745 ;
        RECT  6.640 1.585 6.800 2.425 ;
        RECT  5.925 0.470 6.665 0.630 ;
        RECT  6.585 2.255 6.640 2.425 ;
        RECT  6.425 2.255 6.585 2.495 ;
        RECT  6.250 2.335 6.425 2.495 ;
        RECT  5.805 2.380 5.965 2.540 ;
        RECT  5.805 0.470 5.925 1.715 ;
        RECT  5.765 0.470 5.805 2.540 ;
        RECT  5.125 0.470 5.765 0.630 ;
        RECT  5.645 1.555 5.765 2.540 ;
        RECT  5.455 0.930 5.585 1.375 ;
        RECT  5.425 0.930 5.455 2.540 ;
        RECT  5.295 1.215 5.425 2.540 ;
        RECT  2.855 2.380 5.295 2.540 ;
        RECT  5.025 0.470 5.125 1.020 ;
        RECT  4.965 0.470 5.025 2.165 ;
        RECT  4.865 0.760 4.965 2.165 ;
        RECT  4.655 2.005 4.865 2.165 ;
        RECT  4.405 0.470 4.615 1.195 ;
        RECT  4.245 0.470 4.405 2.200 ;
        RECT  3.235 0.470 4.245 0.785 ;
        RECT  3.165 2.040 4.245 2.200 ;
        RECT  2.915 1.035 3.935 1.295 ;
        RECT  1.595 0.470 3.235 0.630 ;
        RECT  2.655 0.810 2.915 1.295 ;
        RECT  2.695 2.245 2.855 2.540 ;
        RECT  2.275 2.245 2.695 2.405 ;
        RECT  1.935 0.810 2.655 0.970 ;
        RECT  2.355 2.605 2.515 2.880 ;
        RECT  2.275 1.150 2.375 1.310 ;
        RECT  1.935 2.605 2.355 2.765 ;
        RECT  2.115 1.150 2.275 2.405 ;
        RECT  2.015 2.945 2.175 3.220 ;
        RECT  1.595 2.945 2.015 3.105 ;
        RECT  1.775 0.810 1.935 2.765 ;
        RECT  1.435 0.470 1.595 0.755 ;
        RECT  1.435 1.135 1.595 3.105 ;
        RECT  0.385 0.595 1.435 0.755 ;
        RECT  1.425 1.135 1.435 1.295 ;
        RECT  1.295 2.935 1.435 3.105 ;
        RECT  1.165 1.035 1.425 1.295 ;
        RECT  1.035 2.935 1.295 3.195 ;
        RECT  0.895 1.570 1.255 1.830 ;
        RECT  0.635 1.035 0.895 2.555 ;
        RECT  0.385 1.035 0.635 1.195 ;
        RECT  0.125 0.595 0.385 1.195 ;
    END
END ACCSHCINX2

MACRO AFCSIHCONX4
    CLASS CORE ;
    FOREIGN AFCSIHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.635 0.695 10.915 2.895 ;
        END
        ANTENNADIFFAREA     0.7344 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.675 0.595 9.935 0.855 ;
        RECT  9.535 0.595 9.675 0.760 ;
        RECT  9.325 0.470 9.535 0.760 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 0.695 2.255 1.405 ;
        RECT  1.765 2.125 2.025 3.065 ;
        RECT  1.255 1.145 1.965 1.405 ;
        RECT  1.635 2.125 1.765 2.435 ;
        RECT  0.820 2.175 1.635 2.435 ;
        RECT  0.975 0.695 1.255 1.405 ;
        RECT  0.820 1.145 0.975 1.405 ;
        RECT  0.560 1.145 0.820 2.435 ;
        RECT  0.385 1.955 0.560 2.435 ;
        RECT  0.125 1.955 0.385 3.065 ;
        END
        ANTENNADIFFAREA     1.3780 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 2.185 4.065 2.785 ;
        RECT  3.435 2.185 3.805 2.565 ;
        RECT  3.435 0.930 3.680 1.190 ;
        RECT  3.175 0.930 3.435 2.565 ;
        RECT  3.095 2.110 3.175 2.565 ;
        RECT  2.885 2.110 3.095 2.810 ;
        RECT  2.785 2.185 2.885 2.785 ;
        END
        ANTENNADIFFAREA     1.0698 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.145 1.275 4.305 1.665 ;
        RECT  4.050 1.275 4.145 1.435 ;
        RECT  3.890 0.470 4.050 1.435 ;
        RECT  3.805 0.470 3.890 0.760 ;
        RECT  2.905 0.585 3.805 0.745 ;
        RECT  2.745 0.585 2.905 1.745 ;
        RECT  2.645 1.405 2.745 1.745 ;
        RECT  1.375 1.585 2.645 1.745 ;
        RECT  1.115 1.585 1.375 1.845 ;
        END
        ANTENNAGATEAREA     1.2480 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.625 1.595 4.785 2.005 ;
        RECT  4.475 1.845 4.625 2.005 ;
        RECT  4.265 1.845 4.475 2.400 ;
        RECT  3.875 1.845 4.265 2.005 ;
        RECT  3.615 1.715 3.875 2.005 ;
        END
        ANTENNAGATEAREA     1.2077 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.385 -0.250 11.040 0.250 ;
        RECT  10.125 -0.250 10.385 1.075 ;
        RECT  7.655 -0.250 10.125 0.250 ;
        RECT  7.395 -0.250 7.655 0.405 ;
        RECT  6.825 -0.250 7.395 0.250 ;
        RECT  6.665 -0.250 6.825 0.625 ;
        RECT  4.525 -0.250 6.665 0.250 ;
        RECT  4.265 -0.250 4.525 1.095 ;
        RECT  2.825 -0.250 4.265 0.250 ;
        RECT  2.565 -0.250 2.825 0.405 ;
        RECT  1.745 -0.250 2.565 0.250 ;
        RECT  1.485 -0.250 1.745 0.950 ;
        RECT  0.725 -0.250 1.485 0.250 ;
        RECT  0.465 -0.250 0.725 0.945 ;
        RECT  0.000 -0.250 0.465 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.385 3.440 11.040 3.940 ;
        RECT  10.125 2.275 10.385 3.940 ;
        RECT  7.495 3.440 10.125 3.940 ;
        RECT  7.235 3.285 7.495 3.940 ;
        RECT  6.745 3.440 7.235 3.940 ;
        RECT  6.485 3.115 6.745 3.940 ;
        RECT  4.575 3.440 6.485 3.940 ;
        RECT  4.315 2.745 4.575 3.940 ;
        RECT  3.555 3.440 4.315 3.940 ;
        RECT  3.295 2.745 3.555 3.940 ;
        RECT  2.535 3.440 3.295 3.940 ;
        RECT  2.275 2.405 2.535 3.940 ;
        RECT  1.205 3.440 2.275 3.940 ;
        RECT  0.945 2.615 1.205 3.940 ;
        RECT  0.000 3.440 0.945 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.195 1.585 10.455 1.845 ;
        RECT  9.945 1.685 10.195 1.845 ;
        RECT  9.785 1.685 9.945 2.555 ;
        RECT  9.405 2.395 9.785 2.555 ;
        RECT  9.605 1.035 9.735 1.295 ;
        RECT  9.445 1.035 9.605 2.215 ;
        RECT  9.245 1.555 9.445 1.815 ;
        RECT  9.245 2.395 9.405 2.995 ;
        RECT  8.555 2.835 9.245 2.995 ;
        RECT  9.065 1.035 9.225 1.295 ;
        RECT  8.905 0.695 9.065 2.645 ;
        RECT  7.635 0.695 8.905 0.855 ;
        RECT  8.805 2.045 8.905 2.645 ;
        RECT  8.555 1.035 8.715 1.295 ;
        RECT  8.395 1.035 8.555 2.995 ;
        RECT  8.295 2.055 8.395 2.995 ;
        RECT  8.045 1.035 8.205 1.295 ;
        RECT  7.885 1.035 8.045 2.995 ;
        RECT  7.785 2.055 7.885 2.995 ;
        RECT  7.475 0.695 7.635 1.745 ;
        RECT  7.425 1.585 7.475 1.745 ;
        RECT  7.265 1.585 7.425 2.935 ;
        RECT  7.085 0.945 7.295 1.205 ;
        RECT  5.465 2.775 7.265 2.935 ;
        RECT  6.925 0.945 7.085 2.595 ;
        RECT  5.805 2.435 6.925 2.595 ;
        RECT  6.485 1.255 6.585 1.515 ;
        RECT  6.325 0.470 6.485 1.515 ;
        RECT  5.035 0.470 6.325 0.630 ;
        RECT  6.005 1.025 6.145 2.255 ;
        RECT  5.985 0.885 6.005 2.255 ;
        RECT  5.845 0.885 5.985 1.185 ;
        RECT  5.645 1.405 5.805 2.595 ;
        RECT  5.465 0.810 5.545 1.070 ;
        RECT  5.305 0.810 5.465 2.935 ;
        RECT  5.285 0.810 5.305 1.070 ;
        RECT  5.085 1.255 5.125 2.345 ;
        RECT  5.035 1.255 5.085 2.785 ;
        RECT  4.965 0.470 5.035 2.785 ;
        RECT  4.875 0.470 4.965 1.415 ;
        RECT  4.825 2.185 4.965 2.785 ;
        RECT  4.775 0.470 4.875 1.110 ;
    END
END AFCSIHCONX4

MACRO AFCSIHCONX2
    CLASS CORE ;
    FOREIGN AFCSIHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.795 0.695 9.075 2.895 ;
        END
        ANTENNADIFFAREA     0.7344 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.835 0.595 8.095 0.855 ;
        RECT  7.695 0.595 7.835 0.760 ;
        RECT  7.485 0.470 7.695 0.760 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 1.830 1.255 2.895 ;
        RECT  0.335 1.830 0.945 1.990 ;
        RECT  0.715 0.760 0.875 1.135 ;
        RECT  0.335 0.975 0.715 1.135 ;
        RECT  0.125 0.975 0.335 1.990 ;
        END
        ANTENNADIFFAREA     0.6890 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 2.405 2.225 3.005 ;
        RECT  1.715 2.405 1.965 2.565 ;
        RECT  1.595 1.035 1.840 1.295 ;
        RECT  1.595 2.110 1.715 2.565 ;
        RECT  1.555 1.035 1.595 2.565 ;
        RECT  1.505 1.035 1.555 2.400 ;
        RECT  1.435 1.035 1.505 2.335 ;
        END
        ANTENNADIFFAREA     0.6031 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.465 1.405 2.515 1.665 ;
        RECT  2.255 1.255 2.465 1.665 ;
        RECT  2.180 1.255 2.255 1.415 ;
        RECT  2.175 0.600 2.180 1.415 ;
        RECT  2.020 0.470 2.175 1.415 ;
        RECT  1.965 0.470 2.020 0.760 ;
        RECT  1.215 0.590 1.965 0.750 ;
        RECT  1.055 0.590 1.215 1.475 ;
        RECT  0.515 1.315 1.055 1.475 ;
        END
        ANTENNAGATEAREA     0.7631 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.785 1.595 2.945 2.005 ;
        RECT  2.635 1.845 2.785 2.005 ;
        RECT  2.475 1.845 2.635 2.400 ;
        RECT  2.425 2.065 2.475 2.400 ;
        RECT  2.055 2.065 2.425 2.225 ;
        RECT  1.895 1.595 2.055 2.225 ;
        RECT  1.775 1.595 1.895 1.855 ;
        END
        ANTENNAGATEAREA     0.7228 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.545 -0.250 9.200 0.250 ;
        RECT  8.285 -0.250 8.545 1.075 ;
        RECT  5.815 -0.250 8.285 0.250 ;
        RECT  5.555 -0.250 5.815 0.405 ;
        RECT  4.985 -0.250 5.555 0.250 ;
        RECT  4.825 -0.250 4.985 0.625 ;
        RECT  2.685 -0.250 4.825 0.250 ;
        RECT  2.425 -0.250 2.685 1.075 ;
        RECT  1.465 -0.250 2.425 0.250 ;
        RECT  1.205 -0.250 1.465 0.405 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.545 3.440 9.200 3.940 ;
        RECT  8.285 2.275 8.545 3.940 ;
        RECT  5.655 3.440 8.285 3.940 ;
        RECT  5.395 3.285 5.655 3.940 ;
        RECT  4.905 3.440 5.395 3.940 ;
        RECT  4.645 3.115 4.905 3.940 ;
        RECT  2.735 3.440 4.645 3.940 ;
        RECT  2.475 2.640 2.735 3.940 ;
        RECT  1.715 3.440 2.475 3.940 ;
        RECT  1.455 2.745 1.715 3.940 ;
        RECT  0.385 3.440 1.455 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.355 1.585 8.615 1.845 ;
        RECT  8.105 1.685 8.355 1.845 ;
        RECT  7.945 1.685 8.105 2.555 ;
        RECT  7.565 2.395 7.945 2.555 ;
        RECT  7.765 1.035 7.895 1.295 ;
        RECT  7.605 1.035 7.765 2.215 ;
        RECT  7.595 1.555 7.605 2.215 ;
        RECT  7.405 1.555 7.595 1.815 ;
        RECT  7.405 2.395 7.565 2.995 ;
        RECT  6.715 2.835 7.405 2.995 ;
        RECT  7.225 1.035 7.385 1.295 ;
        RECT  7.065 0.695 7.225 2.645 ;
        RECT  5.795 0.695 7.065 0.855 ;
        RECT  6.965 2.045 7.065 2.645 ;
        RECT  6.715 1.035 6.875 1.295 ;
        RECT  6.555 1.035 6.715 2.995 ;
        RECT  6.455 2.055 6.555 2.995 ;
        RECT  6.205 1.035 6.365 1.295 ;
        RECT  6.045 1.035 6.205 2.995 ;
        RECT  5.945 2.055 6.045 2.995 ;
        RECT  5.795 1.585 5.860 1.845 ;
        RECT  5.635 0.695 5.795 1.845 ;
        RECT  5.585 1.685 5.635 1.845 ;
        RECT  5.425 1.685 5.585 2.935 ;
        RECT  5.245 0.945 5.455 1.205 ;
        RECT  3.625 2.775 5.425 2.935 ;
        RECT  5.085 0.945 5.245 2.595 ;
        RECT  3.965 2.435 5.085 2.595 ;
        RECT  4.645 1.255 4.745 1.515 ;
        RECT  4.485 0.470 4.645 1.515 ;
        RECT  3.195 0.470 4.485 0.630 ;
        RECT  4.145 0.885 4.305 2.255 ;
        RECT  3.955 0.885 4.145 1.145 ;
        RECT  3.805 1.405 3.965 2.595 ;
        RECT  3.625 0.810 3.705 1.070 ;
        RECT  3.465 0.810 3.625 2.935 ;
        RECT  3.445 0.810 3.465 1.070 ;
        RECT  3.245 1.255 3.285 2.345 ;
        RECT  3.195 1.255 3.245 2.785 ;
        RECT  3.125 0.470 3.195 2.785 ;
        RECT  3.035 0.470 3.125 1.415 ;
        RECT  2.985 2.185 3.125 2.785 ;
        RECT  2.935 0.470 3.035 1.110 ;
    END
END AFCSIHCONX2

MACRO AFCSHCONX4
    CLASS CORE ;
    FOREIGN AFCSHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  27.475 0.595 27.495 2.585 ;
        RECT  27.265 0.595 27.475 3.045 ;
        RECT  27.215 2.105 27.265 3.045 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  26.805 0.880 27.015 1.170 ;
        RECT  26.695 1.010 26.805 1.170 ;
        RECT  26.535 1.010 26.695 1.755 ;
        RECT  26.365 1.495 26.535 1.755 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.435 1.545 18.900 1.705 ;
        RECT  16.435 2.565 18.900 2.725 ;
        RECT  16.250 1.545 16.435 2.725 ;
        RECT  16.225 1.700 16.250 2.520 ;
        END
        ANTENNADIFFAREA     1.8708 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.760 2.605 16.020 2.865 ;
        RECT  14.970 2.655 15.760 2.815 ;
        RECT  14.710 2.605 14.970 2.865 ;
        RECT  14.410 2.605 14.710 2.815 ;
        RECT  14.255 1.490 14.590 1.650 ;
        RECT  14.255 2.520 14.410 2.815 ;
        RECT  14.230 1.490 14.255 2.815 ;
        RECT  13.970 1.490 14.230 2.860 ;
        RECT  13.950 1.490 13.970 2.810 ;
        RECT  13.250 1.490 13.950 1.750 ;
        RECT  13.925 1.990 13.950 2.810 ;
        RECT  13.215 2.325 13.925 2.485 ;
        RECT  13.210 2.325 13.215 2.585 ;
        RECT  13.050 2.325 13.210 2.860 ;
        RECT  12.950 2.600 13.050 2.860 ;
        END
        ANTENNADIFFAREA     1.6968 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.415 1.715 22.430 1.975 ;
        RECT  22.205 1.700 22.415 1.990 ;
        RECT  21.490 1.715 22.205 1.975 ;
        END
        ANTENNAGATEAREA     0.9516 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.780 7.695 2.040 ;
        RECT  6.755 1.780 6.775 2.400 ;
        RECT  6.615 1.880 6.755 2.400 ;
        RECT  6.565 2.110 6.615 2.400 ;
        END
        ANTENNAGATEAREA     0.9516 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.635 4.475 1.990 ;
        RECT  3.955 1.635 4.265 1.850 ;
        END
        ANTENNAGATEAREA     0.7735 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.555 0.875 1.990 ;
        RECT  0.515 1.555 0.585 1.815 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.935 -0.250 27.600 0.250 ;
        RECT  26.675 -0.250 26.935 0.405 ;
        RECT  25.670 -0.250 26.675 0.250 ;
        RECT  25.410 -0.250 25.670 0.575 ;
        RECT  23.570 -0.250 25.410 0.250 ;
        RECT  23.310 -0.250 23.570 0.405 ;
        RECT  22.430 -0.250 23.310 0.250 ;
        RECT  22.170 -0.250 22.430 0.405 ;
        RECT  21.270 -0.250 22.170 0.250 ;
        RECT  21.010 -0.250 21.270 0.405 ;
        RECT  9.600 -0.250 21.010 0.250 ;
        RECT  9.440 -0.250 9.600 1.235 ;
        RECT  7.510 -0.250 9.440 0.250 ;
        RECT  6.570 -0.250 7.510 0.575 ;
        RECT  5.300 -0.250 6.570 0.250 ;
        RECT  5.040 -0.250 5.300 0.405 ;
        RECT  4.430 -0.250 5.040 0.250 ;
        RECT  4.170 -0.250 4.430 0.405 ;
        RECT  1.810 -0.250 4.170 0.250 ;
        RECT  1.550 -0.250 1.810 0.405 ;
        RECT  0.895 -0.250 1.550 0.250 ;
        RECT  0.635 -0.250 0.895 1.195 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.935 3.440 27.600 3.940 ;
        RECT  26.675 2.825 26.935 3.940 ;
        RECT  26.350 3.440 26.675 3.940 ;
        RECT  26.090 2.745 26.350 3.940 ;
        RECT  23.520 3.440 26.090 3.940 ;
        RECT  23.260 2.415 23.520 3.940 ;
        RECT  22.470 3.405 23.260 3.940 ;
        RECT  22.210 3.285 22.470 3.940 ;
        RECT  21.390 3.440 22.210 3.940 ;
        RECT  21.130 3.285 21.390 3.940 ;
        RECT  10.500 3.440 21.130 3.940 ;
        RECT  10.240 3.115 10.500 3.940 ;
        RECT  9.865 3.440 10.240 3.940 ;
        RECT  9.605 3.285 9.865 3.940 ;
        RECT  8.775 3.440 9.605 3.940 ;
        RECT  8.515 3.285 8.775 3.940 ;
        RECT  7.725 3.440 8.515 3.940 ;
        RECT  7.465 3.125 7.725 3.940 ;
        RECT  6.635 3.440 7.465 3.940 ;
        RECT  6.375 3.285 6.635 3.940 ;
        RECT  5.685 3.440 6.375 3.940 ;
        RECT  5.425 3.285 5.685 3.940 ;
        RECT  4.530 3.440 5.425 3.940 ;
        RECT  4.270 3.285 4.530 3.940 ;
        RECT  1.805 3.440 4.270 3.940 ;
        RECT  1.545 2.945 1.805 3.940 ;
        RECT  0.895 3.440 1.545 3.940 ;
        RECT  0.635 2.935 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  27.035 1.495 27.055 1.755 ;
        RECT  26.875 1.495 27.035 2.565 ;
        RECT  25.890 2.405 26.875 2.565 ;
        RECT  26.155 2.065 26.395 2.225 ;
        RECT  26.155 1.035 26.355 1.295 ;
        RECT  25.995 1.035 26.155 2.225 ;
        RECT  25.550 2.065 25.995 2.225 ;
        RECT  25.730 2.405 25.890 3.220 ;
        RECT  24.530 3.060 25.730 3.220 ;
        RECT  25.645 1.425 25.695 1.685 ;
        RECT  25.485 0.755 25.645 1.685 ;
        RECT  25.390 2.065 25.550 2.880 ;
        RECT  25.105 0.755 25.485 0.915 ;
        RECT  25.435 1.425 25.485 1.685 ;
        RECT  24.870 2.720 25.390 2.880 ;
        RECT  25.050 1.095 25.210 2.540 ;
        RECT  24.945 0.585 25.105 0.915 ;
        RECT  24.870 1.095 25.050 1.255 ;
        RECT  19.360 0.585 24.945 0.745 ;
        RECT  24.710 1.445 24.870 2.880 ;
        RECT  24.450 0.925 24.620 1.185 ;
        RECT  24.450 2.320 24.530 3.220 ;
        RECT  24.370 0.925 24.450 3.220 ;
        RECT  24.290 0.925 24.370 2.485 ;
        RECT  23.850 0.925 24.110 3.090 ;
        RECT  23.810 2.150 23.850 3.090 ;
        RECT  23.510 0.925 23.670 1.660 ;
        RECT  20.360 0.925 23.510 1.085 ;
        RECT  22.950 2.165 23.010 3.105 ;
        RECT  22.950 1.265 23.000 1.425 ;
        RECT  22.790 1.265 22.950 3.105 ;
        RECT  22.740 1.265 22.790 1.425 ;
        RECT  22.750 2.165 22.790 3.105 ;
        RECT  19.345 2.945 22.750 3.105 ;
        RECT  21.670 2.165 21.930 2.765 ;
        RECT  21.310 1.265 21.850 1.425 ;
        RECT  21.310 2.165 21.670 2.325 ;
        RECT  19.930 2.605 21.670 2.765 ;
        RECT  21.150 1.265 21.310 2.325 ;
        RECT  20.950 1.725 21.150 1.985 ;
        RECT  20.770 2.165 20.950 2.425 ;
        RECT  20.770 1.265 20.800 1.425 ;
        RECT  20.610 1.265 20.770 2.425 ;
        RECT  20.540 1.265 20.610 1.425 ;
        RECT  20.360 2.165 20.390 2.425 ;
        RECT  20.200 0.925 20.360 2.425 ;
        RECT  20.000 0.925 20.200 1.185 ;
        RECT  19.700 2.165 19.930 2.765 ;
        RECT  19.540 0.935 19.700 2.765 ;
        RECT  19.200 0.585 19.360 1.365 ;
        RECT  19.185 2.055 19.345 3.105 ;
        RECT  15.875 1.205 19.200 1.365 ;
        RECT  18.900 2.055 19.185 2.215 ;
        RECT  18.860 0.525 19.020 0.785 ;
        RECT  18.300 2.005 18.900 2.265 ;
        RECT  15.890 0.525 18.860 0.685 ;
        RECT  15.710 0.865 18.620 1.025 ;
        RECT  17.325 2.055 18.300 2.215 ;
        RECT  17.775 2.905 17.825 3.165 ;
        RECT  17.565 2.905 17.775 3.220 ;
        RECT  14.340 3.060 17.565 3.220 ;
        RECT  16.725 2.005 17.325 2.265 ;
        RECT  15.715 1.205 15.875 2.415 ;
        RECT  14.935 2.255 15.715 2.415 ;
        RECT  15.550 0.470 15.710 1.025 ;
        RECT  9.940 0.470 15.550 0.630 ;
        RECT  15.370 1.475 15.510 2.075 ;
        RECT  15.210 0.810 15.370 2.075 ;
        RECT  10.280 0.810 15.210 0.970 ;
        RECT  14.775 1.150 14.935 2.415 ;
        RECT  11.520 1.150 14.775 1.310 ;
        RECT  13.620 2.670 13.720 2.930 ;
        RECT  13.460 2.670 13.620 3.220 ;
        RECT  12.700 3.060 13.460 3.220 ;
        RECT  12.790 1.490 12.950 2.045 ;
        RECT  12.650 1.885 12.790 2.045 ;
        RECT  12.650 2.720 12.700 3.220 ;
        RECT  12.490 1.885 12.650 3.220 ;
        RECT  12.080 1.490 12.490 1.650 ;
        RECT  12.440 2.720 12.490 3.220 ;
        RECT  10.840 3.060 12.440 3.220 ;
        RECT  12.080 2.620 12.110 2.880 ;
        RECT  11.920 1.490 12.080 2.880 ;
        RECT  11.850 2.620 11.920 2.880 ;
        RECT  11.180 2.720 11.850 2.880 ;
        RECT  11.360 1.150 11.520 2.540 ;
        RECT  11.310 1.150 11.360 1.310 ;
        RECT  11.020 2.435 11.180 2.880 ;
        RECT  11.010 1.150 11.060 1.310 ;
        RECT  11.010 2.095 11.060 2.255 ;
        RECT  10.620 2.435 11.020 2.595 ;
        RECT  10.850 1.150 11.010 2.255 ;
        RECT  10.800 1.150 10.850 1.310 ;
        RECT  10.800 2.095 10.850 2.255 ;
        RECT  10.680 2.775 10.840 3.220 ;
        RECT  10.060 2.775 10.680 2.935 ;
        RECT  10.460 1.675 10.620 2.595 ;
        RECT  9.705 2.435 10.460 2.595 ;
        RECT  10.120 0.810 10.280 2.255 ;
        RECT  9.325 2.095 10.120 2.255 ;
        RECT  9.900 2.775 10.060 3.105 ;
        RECT  9.780 0.470 9.940 1.915 ;
        RECT  8.415 2.945 9.900 3.105 ;
        RECT  8.920 1.755 9.780 1.915 ;
        RECT  9.545 2.435 9.705 2.765 ;
        RECT  9.260 1.415 9.600 1.575 ;
        RECT  8.755 2.605 9.545 2.765 ;
        RECT  9.065 2.095 9.325 2.425 ;
        RECT  9.100 0.470 9.260 1.575 ;
        RECT  7.900 0.470 9.100 0.630 ;
        RECT  8.580 2.095 9.065 2.255 ;
        RECT  8.760 0.810 8.920 1.915 ;
        RECT  8.240 0.810 8.760 0.970 ;
        RECT  8.595 2.445 8.755 2.765 ;
        RECT  8.215 2.445 8.595 2.605 ;
        RECT  8.420 1.150 8.580 2.255 ;
        RECT  8.255 2.785 8.415 3.105 ;
        RECT  6.775 2.785 8.255 2.945 ;
        RECT  8.080 0.810 8.240 1.255 ;
        RECT  8.055 1.435 8.215 2.605 ;
        RECT  6.230 1.095 8.080 1.255 ;
        RECT  6.530 1.435 8.055 1.595 ;
        RECT  7.135 2.445 8.055 2.605 ;
        RECT  7.740 0.470 7.900 0.915 ;
        RECT  5.850 0.755 7.740 0.915 ;
        RECT  6.975 2.320 7.135 2.605 ;
        RECT  6.615 2.785 6.775 3.105 ;
        RECT  4.095 2.945 6.615 3.105 ;
        RECT  6.135 2.605 6.235 2.765 ;
        RECT  6.070 1.095 6.230 2.085 ;
        RECT  5.975 2.265 6.135 2.765 ;
        RECT  5.155 1.925 6.070 2.085 ;
        RECT  4.815 2.265 5.975 2.425 ;
        RECT  5.750 0.755 5.850 1.155 ;
        RECT  5.590 0.610 5.750 1.155 ;
        RECT  4.350 0.610 5.590 0.770 ;
        RECT  2.855 2.605 5.465 2.765 ;
        RECT  4.995 0.950 5.155 2.085 ;
        RECT  4.640 0.950 4.995 1.110 ;
        RECT  4.655 1.290 4.815 2.425 ;
        RECT  4.350 1.290 4.655 1.450 ;
        RECT  4.190 0.610 4.350 1.450 ;
        RECT  3.935 2.945 4.095 3.140 ;
        RECT  2.240 2.980 3.935 3.140 ;
        RECT  3.720 0.685 3.890 1.285 ;
        RECT  3.720 2.145 3.875 2.405 ;
        RECT  3.630 0.685 3.720 2.405 ;
        RECT  3.560 1.125 3.630 2.405 ;
        RECT  3.390 1.605 3.560 1.865 ;
        RECT  3.210 0.705 3.380 1.305 ;
        RECT  3.210 2.165 3.365 2.425 ;
        RECT  3.050 0.585 3.210 2.425 ;
        RECT  1.405 0.585 3.050 0.745 ;
        RECT  2.770 0.965 2.870 1.125 ;
        RECT  2.770 2.200 2.855 2.800 ;
        RECT  2.610 0.965 2.770 2.800 ;
        RECT  2.595 2.200 2.610 2.800 ;
        RECT  2.260 0.965 2.360 1.125 ;
        RECT  2.260 2.155 2.345 2.415 ;
        RECT  2.100 0.965 2.260 2.415 ;
        RECT  2.080 2.595 2.240 3.140 ;
        RECT  2.085 2.155 2.100 2.415 ;
        RECT  0.385 2.595 2.080 2.755 ;
        RECT  1.405 1.550 1.780 1.810 ;
        RECT  1.245 0.585 1.405 2.300 ;
        RECT  1.145 1.035 1.245 1.295 ;
        RECT  1.145 2.040 1.245 2.300 ;
        RECT  0.335 0.695 0.385 1.295 ;
        RECT  0.335 2.105 0.385 3.045 ;
        RECT  0.175 0.695 0.335 3.045 ;
        RECT  0.125 0.695 0.175 1.295 ;
        RECT  0.125 2.105 0.175 3.045 ;
    END
END AFCSHCONX4

MACRO AFCSHCONX2
    CLASS CORE ;
    FOREIGN AFCSHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 23.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.795 0.595 23.815 2.585 ;
        RECT  23.585 0.595 23.795 3.045 ;
        RECT  23.535 2.105 23.585 3.045 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.125 0.880 23.335 1.170 ;
        RECT  23.015 1.010 23.125 1.170 ;
        RECT  22.855 1.010 23.015 1.755 ;
        RECT  22.685 1.495 22.855 1.755 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.410 1.700 16.435 2.400 ;
        RECT  16.225 1.630 16.410 2.400 ;
        RECT  13.730 1.630 16.225 1.790 ;
        RECT  13.905 2.630 14.515 2.890 ;
        RECT  13.730 2.630 13.905 2.790 ;
        RECT  13.570 1.630 13.730 2.790 ;
        RECT  13.480 1.630 13.570 1.790 ;
        END
        ANTENNADIFFAREA     1.3509 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.220 3.060 13.520 3.220 ;
        RECT  12.060 2.240 12.220 3.220 ;
        RECT  11.835 2.240 12.060 2.400 ;
        RECT  11.835 1.490 11.985 1.650 ;
        RECT  11.650 1.490 11.835 2.400 ;
        RECT  11.625 1.700 11.650 2.400 ;
        RECT  11.200 2.240 11.625 2.400 ;
        RECT  11.040 2.240 11.200 2.830 ;
        END
        ANTENNADIFFAREA     1.1994 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.735 1.715 19.060 1.975 ;
        RECT  18.525 1.700 18.735 1.990 ;
        RECT  18.460 1.715 18.525 1.975 ;
        END
        ANTENNAGATEAREA     0.4758 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 1.790 7.260 2.050 ;
        RECT  7.025 1.790 7.235 2.400 ;
        RECT  7.000 1.790 7.025 2.050 ;
        END
        ANTENNAGATEAREA     0.4784 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.635 4.475 1.990 ;
        RECT  3.955 1.635 4.265 1.850 ;
        END
        ANTENNAGATEAREA     0.7735 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.555 0.875 1.990 ;
        RECT  0.515 1.555 0.585 1.815 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  23.255 -0.250 23.920 0.250 ;
        RECT  22.995 -0.250 23.255 0.405 ;
        RECT  21.990 -0.250 22.995 0.250 ;
        RECT  21.730 -0.250 21.990 0.575 ;
        RECT  19.890 -0.250 21.730 0.250 ;
        RECT  19.630 -0.250 19.890 0.405 ;
        RECT  18.260 -0.250 19.630 0.250 ;
        RECT  18.000 -0.250 18.260 0.405 ;
        RECT  8.690 -0.250 18.000 0.250 ;
        RECT  8.090 -0.250 8.690 0.575 ;
        RECT  7.260 -0.250 8.090 0.250 ;
        RECT  6.320 -0.250 7.260 0.575 ;
        RECT  5.300 -0.250 6.320 0.250 ;
        RECT  5.040 -0.250 5.300 0.405 ;
        RECT  4.430 -0.250 5.040 0.250 ;
        RECT  4.170 -0.250 4.430 0.405 ;
        RECT  1.810 -0.250 4.170 0.250 ;
        RECT  1.550 -0.250 1.810 0.405 ;
        RECT  0.895 -0.250 1.550 0.250 ;
        RECT  0.635 -0.250 0.895 1.195 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  23.255 3.440 23.920 3.940 ;
        RECT  22.995 2.825 23.255 3.940 ;
        RECT  22.670 3.440 22.995 3.940 ;
        RECT  22.410 2.745 22.670 3.940 ;
        RECT  19.900 3.440 22.410 3.940 ;
        RECT  19.640 2.150 19.900 3.940 ;
        RECT  18.340 3.440 19.640 3.940 ;
        RECT  18.080 3.285 18.340 3.940 ;
        RECT  8.915 3.440 18.080 3.940 ;
        RECT  8.655 3.115 8.915 3.940 ;
        RECT  7.725 3.440 8.655 3.940 ;
        RECT  7.465 3.285 7.725 3.940 ;
        RECT  6.635 3.440 7.465 3.940 ;
        RECT  6.375 3.285 6.635 3.940 ;
        RECT  5.685 3.440 6.375 3.940 ;
        RECT  5.425 3.285 5.685 3.940 ;
        RECT  4.530 3.440 5.425 3.940 ;
        RECT  4.270 3.285 4.530 3.940 ;
        RECT  1.805 3.440 4.270 3.940 ;
        RECT  1.545 2.945 1.805 3.940 ;
        RECT  0.895 3.440 1.545 3.940 ;
        RECT  0.635 2.935 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  23.355 1.495 23.375 1.755 ;
        RECT  23.195 1.495 23.355 2.565 ;
        RECT  22.230 2.405 23.195 2.565 ;
        RECT  22.475 2.065 22.715 2.225 ;
        RECT  22.475 1.035 22.675 1.295 ;
        RECT  22.315 1.035 22.475 2.225 ;
        RECT  21.890 2.065 22.315 2.225 ;
        RECT  22.070 2.405 22.230 3.220 ;
        RECT  20.870 3.060 22.070 3.220 ;
        RECT  21.965 1.425 22.015 1.685 ;
        RECT  21.805 0.755 21.965 1.685 ;
        RECT  21.730 2.065 21.890 2.880 ;
        RECT  21.365 0.755 21.805 0.915 ;
        RECT  21.755 1.425 21.805 1.685 ;
        RECT  21.210 2.720 21.730 2.880 ;
        RECT  21.390 1.095 21.550 2.540 ;
        RECT  21.190 1.095 21.390 1.255 ;
        RECT  21.205 0.585 21.365 0.915 ;
        RECT  21.050 1.445 21.210 2.880 ;
        RECT  16.350 0.585 21.205 0.745 ;
        RECT  20.870 0.925 20.940 1.185 ;
        RECT  20.710 0.925 20.870 3.220 ;
        RECT  20.680 0.925 20.710 1.185 ;
        RECT  20.170 0.925 20.430 3.090 ;
        RECT  20.150 2.150 20.170 3.090 ;
        RECT  19.830 0.925 19.990 1.845 ;
        RECT  17.350 0.925 19.830 1.085 ;
        RECT  19.240 1.265 19.400 3.105 ;
        RECT  19.090 1.265 19.240 1.425 ;
        RECT  19.130 2.165 19.240 3.105 ;
        RECT  15.890 2.945 19.130 3.105 ;
        RECT  18.620 2.170 18.880 2.765 ;
        RECT  18.280 1.265 18.800 1.425 ;
        RECT  18.280 2.170 18.620 2.330 ;
        RECT  16.920 2.605 18.620 2.765 ;
        RECT  18.120 1.265 18.280 2.330 ;
        RECT  17.940 1.725 18.120 1.985 ;
        RECT  17.760 2.165 17.940 2.425 ;
        RECT  17.760 1.265 17.790 1.425 ;
        RECT  17.600 1.265 17.760 2.425 ;
        RECT  17.530 1.265 17.600 1.425 ;
        RECT  17.350 2.165 17.380 2.425 ;
        RECT  17.190 0.925 17.350 2.425 ;
        RECT  16.990 0.925 17.190 1.185 ;
        RECT  16.775 2.165 16.920 2.765 ;
        RECT  16.615 0.935 16.775 2.765 ;
        RECT  16.530 0.935 16.615 1.195 ;
        RECT  16.190 0.585 16.350 1.450 ;
        RECT  13.300 1.290 16.190 1.450 ;
        RECT  13.420 0.580 16.010 0.740 ;
        RECT  13.240 0.950 15.890 1.110 ;
        RECT  15.730 2.090 15.890 3.105 ;
        RECT  15.290 2.090 15.730 2.350 ;
        RECT  14.510 2.170 15.290 2.330 ;
        RECT  13.910 2.120 14.510 2.380 ;
        RECT  13.140 1.290 13.300 2.880 ;
        RECT  13.080 0.470 13.240 1.110 ;
        RECT  12.560 2.720 13.140 2.880 ;
        RECT  9.030 0.470 13.080 0.630 ;
        RECT  12.740 0.810 12.900 2.540 ;
        RECT  9.370 0.810 12.740 0.970 ;
        RECT  12.400 1.150 12.560 2.880 ;
        RECT  10.150 1.150 12.400 1.310 ;
        RECT  11.660 2.580 11.760 2.840 ;
        RECT  11.500 2.580 11.660 3.220 ;
        RECT  10.860 3.060 11.500 3.220 ;
        RECT  11.245 1.490 11.415 1.650 ;
        RECT  11.085 1.490 11.245 2.010 ;
        RECT  10.860 1.850 11.085 2.010 ;
        RECT  10.520 1.490 10.905 1.650 ;
        RECT  10.700 1.850 10.860 3.220 ;
        RECT  9.710 3.060 10.700 3.220 ;
        RECT  10.360 1.490 10.520 2.860 ;
        RECT  10.265 2.435 10.360 2.860 ;
        RECT  9.035 2.435 10.265 2.595 ;
        RECT  9.990 1.150 10.150 2.255 ;
        RECT  9.725 2.095 9.990 2.255 ;
        RECT  9.710 1.150 9.810 1.310 ;
        RECT  9.550 1.150 9.710 1.725 ;
        RECT  9.550 2.775 9.710 3.220 ;
        RECT  9.480 1.565 9.550 1.725 ;
        RECT  8.275 2.775 9.550 2.935 ;
        RECT  9.320 1.565 9.480 2.255 ;
        RECT  9.210 0.810 9.370 1.255 ;
        RECT  9.215 2.095 9.320 2.255 ;
        RECT  8.695 1.095 9.210 1.255 ;
        RECT  8.875 1.675 9.035 2.595 ;
        RECT  8.870 0.470 9.030 0.915 ;
        RECT  7.720 2.435 8.875 2.595 ;
        RECT  6.140 0.755 8.870 0.915 ;
        RECT  8.535 1.095 8.695 2.255 ;
        RECT  7.630 1.095 8.535 1.255 ;
        RECT  8.035 2.095 8.535 2.255 ;
        RECT  8.195 1.435 8.355 1.915 ;
        RECT  8.115 2.775 8.275 3.105 ;
        RECT  7.325 1.435 8.195 1.595 ;
        RECT  2.150 2.945 8.115 3.105 ;
        RECT  7.560 2.435 7.720 2.740 ;
        RECT  6.820 2.580 7.560 2.740 ;
        RECT  7.165 1.095 7.325 1.595 ;
        RECT  6.480 1.095 7.165 1.255 ;
        RECT  6.820 1.435 6.920 1.595 ;
        RECT  6.660 1.435 6.820 2.740 ;
        RECT  6.320 1.095 6.480 2.425 ;
        RECT  6.235 2.265 6.320 2.425 ;
        RECT  5.975 2.265 6.235 2.745 ;
        RECT  5.980 0.755 6.140 2.085 ;
        RECT  5.155 1.925 5.980 2.085 ;
        RECT  4.815 2.265 5.975 2.425 ;
        RECT  5.640 0.610 5.800 1.095 ;
        RECT  4.350 0.610 5.640 0.770 ;
        RECT  2.855 2.605 5.465 2.765 ;
        RECT  4.995 0.950 5.155 2.085 ;
        RECT  4.640 0.950 4.995 1.110 ;
        RECT  4.655 1.290 4.815 2.425 ;
        RECT  4.350 1.290 4.655 1.450 ;
        RECT  4.190 0.610 4.350 1.450 ;
        RECT  3.720 0.685 3.890 1.285 ;
        RECT  3.720 2.145 3.875 2.405 ;
        RECT  3.630 0.685 3.720 2.405 ;
        RECT  3.560 1.125 3.630 2.405 ;
        RECT  3.390 1.605 3.560 1.865 ;
        RECT  3.210 0.705 3.380 1.305 ;
        RECT  3.210 2.165 3.365 2.425 ;
        RECT  3.050 0.585 3.210 2.425 ;
        RECT  1.405 0.585 3.050 0.745 ;
        RECT  2.770 0.965 2.870 1.125 ;
        RECT  2.770 2.165 2.855 2.765 ;
        RECT  2.610 0.965 2.770 2.765 ;
        RECT  2.595 2.165 2.610 2.765 ;
        RECT  2.260 0.965 2.360 1.125 ;
        RECT  2.260 2.155 2.345 2.415 ;
        RECT  2.100 0.965 2.260 2.415 ;
        RECT  1.990 2.595 2.150 3.105 ;
        RECT  2.085 2.155 2.100 2.415 ;
        RECT  0.385 2.595 1.990 2.755 ;
        RECT  1.405 1.550 1.780 1.810 ;
        RECT  1.245 0.585 1.405 2.300 ;
        RECT  1.145 1.035 1.245 1.295 ;
        RECT  1.145 2.040 1.245 2.300 ;
        RECT  0.335 0.695 0.385 1.295 ;
        RECT  0.335 2.105 0.385 3.045 ;
        RECT  0.175 0.695 0.335 3.045 ;
        RECT  0.125 0.695 0.175 1.295 ;
        RECT  0.125 2.105 0.175 3.045 ;
    END
END AFCSHCONX2

MACRO AFCSHCINX4
    CLASS CORE ;
    FOREIGN AFCSHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  27.015 0.595 27.020 2.335 ;
        RECT  26.995 0.595 27.015 2.995 ;
        RECT  26.805 0.595 26.995 3.195 ;
        RECT  26.735 0.595 26.805 1.195 ;
        RECT  26.735 2.255 26.805 3.195 ;
        END
        ANTENNADIFFAREA     0.7250 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  26.345 0.880 26.555 1.170 ;
        RECT  26.085 1.010 26.345 1.170 ;
        RECT  25.925 1.010 26.085 1.755 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.975 1.610 18.490 1.870 ;
        RECT  15.975 2.630 18.400 2.890 ;
        RECT  15.765 1.610 15.975 2.890 ;
        RECT  15.750 1.610 15.765 1.870 ;
        RECT  15.750 2.630 15.765 2.890 ;
        END
        ANTENNADIFFAREA     1.5552 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.055 2.460 15.065 2.720 ;
        RECT  14.845 1.490 15.055 2.810 ;
        RECT  14.005 1.490 14.845 1.720 ;
        RECT  14.125 2.460 14.845 2.720 ;
        RECT  14.110 2.540 14.125 2.720 ;
        RECT  13.030 2.540 14.110 2.700 ;
        RECT  13.015 1.490 14.005 1.650 ;
        RECT  12.415 2.540 13.030 2.800 ;
        RECT  12.415 1.490 13.015 1.750 ;
        END
        ANTENNADIFFAREA     1.8708 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.125 1.700 22.640 1.990 ;
        END
        ANTENNAGATEAREA     0.5590 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.415 1.565 7.720 2.075 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.055 1.605 7.235 2.000 ;
        RECT  6.895 1.605 7.055 2.420 ;
        RECT  6.800 1.605 6.895 2.000 ;
        RECT  5.250 2.260 6.895 2.420 ;
        RECT  6.725 1.605 6.800 1.765 ;
        RECT  5.215 2.255 5.250 2.515 ;
        RECT  5.055 1.770 5.215 2.515 ;
        RECT  5.050 1.770 5.055 1.930 ;
        RECT  4.890 0.925 5.050 1.930 ;
        END
        ANTENNAGATEAREA     0.6864 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.495 0.915 1.990 ;
        RECT  0.465 1.495 0.585 1.755 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.325 -0.250 27.140 0.250 ;
        RECT  26.065 -0.250 26.325 0.405 ;
        RECT  25.465 -0.250 26.065 0.250 ;
        RECT  25.205 -0.250 25.465 0.785 ;
        RECT  23.115 -0.250 25.205 0.250 ;
        RECT  22.855 -0.250 23.115 0.405 ;
        RECT  21.830 -0.250 22.855 0.250 ;
        RECT  20.890 -0.250 21.830 0.405 ;
        RECT  6.030 -0.250 20.890 0.250 ;
        RECT  5.770 -0.250 6.030 0.405 ;
        RECT  1.865 -0.250 5.770 0.250 ;
        RECT  1.605 -0.250 1.865 0.405 ;
        RECT  0.925 -0.250 1.605 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.435 3.440 27.140 3.940 ;
        RECT  26.175 2.800 26.435 3.940 ;
        RECT  25.775 3.440 26.175 3.940 ;
        RECT  25.515 2.745 25.775 3.940 ;
        RECT  23.005 3.440 25.515 3.940 ;
        RECT  22.745 2.165 23.005 3.940 ;
        RECT  21.780 3.440 22.745 3.940 ;
        RECT  20.840 3.285 21.780 3.940 ;
        RECT  7.950 3.440 20.840 3.940 ;
        RECT  7.010 3.285 7.950 3.940 ;
        RECT  1.805 3.440 7.010 3.940 ;
        RECT  1.545 3.285 1.805 3.940 ;
        RECT  0.895 3.440 1.545 3.940 ;
        RECT  0.635 2.255 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  26.445 1.495 26.605 2.055 ;
        RECT  26.430 1.895 26.445 2.055 ;
        RECT  26.270 1.895 26.430 2.565 ;
        RECT  25.335 2.405 26.270 2.565 ;
        RECT  25.695 1.965 25.895 2.225 ;
        RECT  25.695 1.035 25.745 1.295 ;
        RECT  25.535 1.035 25.695 2.225 ;
        RECT  25.485 1.035 25.535 1.295 ;
        RECT  24.995 2.065 25.535 2.225 ;
        RECT  25.175 2.405 25.335 3.220 ;
        RECT  23.975 3.060 25.175 3.220 ;
        RECT  25.020 1.465 25.120 1.725 ;
        RECT  24.860 0.585 25.020 1.725 ;
        RECT  24.835 2.065 24.995 2.880 ;
        RECT  19.080 0.585 24.860 0.745 ;
        RECT  24.315 2.720 24.835 2.880 ;
        RECT  24.655 1.005 24.680 1.265 ;
        RECT  24.495 1.005 24.655 2.540 ;
        RECT  24.420 1.005 24.495 1.265 ;
        RECT  24.155 1.445 24.315 2.880 ;
        RECT  23.975 0.925 24.170 1.185 ;
        RECT  23.815 0.925 23.975 3.220 ;
        RECT  23.525 0.925 23.610 1.185 ;
        RECT  23.515 0.925 23.525 2.700 ;
        RECT  23.365 0.925 23.515 3.090 ;
        RECT  23.255 2.150 23.365 3.090 ;
        RECT  23.045 1.645 23.175 1.905 ;
        RECT  22.885 0.925 23.045 1.905 ;
        RECT  20.030 0.925 22.885 1.085 ;
        RECT  21.945 1.265 22.545 1.425 ;
        RECT  22.235 2.195 22.495 3.135 ;
        RECT  21.945 2.585 22.235 2.880 ;
        RECT  21.785 1.265 21.945 2.880 ;
        RECT  19.540 2.720 21.785 2.880 ;
        RECT  21.500 1.265 21.595 1.425 ;
        RECT  21.340 1.265 21.500 2.500 ;
        RECT  21.335 1.265 21.340 1.970 ;
        RECT  20.900 1.810 21.335 1.970 ;
        RECT  20.640 1.760 20.900 2.020 ;
        RECT  20.460 1.265 20.570 1.425 ;
        RECT  20.460 2.245 20.560 2.505 ;
        RECT  20.300 1.265 20.460 2.505 ;
        RECT  19.980 2.245 20.050 2.505 ;
        RECT  19.980 0.925 20.030 1.185 ;
        RECT  19.820 0.925 19.980 2.505 ;
        RECT  19.770 0.925 19.820 1.185 ;
        RECT  19.790 2.245 19.820 2.505 ;
        RECT  19.280 0.925 19.540 2.880 ;
        RECT  19.260 0.925 19.280 1.185 ;
        RECT  16.420 2.120 19.280 2.380 ;
        RECT  18.920 0.585 19.080 1.160 ;
        RECT  18.400 1.000 18.920 1.160 ;
        RECT  18.580 0.470 18.740 0.820 ;
        RECT  6.370 0.470 18.580 0.630 ;
        RECT  18.240 0.810 18.400 1.160 ;
        RECT  15.020 0.810 18.240 0.970 ;
        RECT  15.540 1.150 18.060 1.310 ;
        RECT  15.380 1.150 15.540 3.220 ;
        RECT  8.920 3.060 15.380 3.220 ;
        RECT  14.860 0.810 15.020 1.310 ;
        RECT  10.910 1.150 14.860 1.310 ;
        RECT  6.710 0.810 14.600 0.970 ;
        RECT  14.000 1.950 14.600 2.240 ;
        RECT  13.015 2.080 14.000 2.240 ;
        RECT  12.415 2.030 13.015 2.290 ;
        RECT  12.020 2.080 12.415 2.240 ;
        RECT  12.020 1.495 12.025 1.655 ;
        RECT  11.860 1.495 12.020 2.880 ;
        RECT  11.765 1.495 11.860 1.655 ;
        RECT  10.120 2.720 11.860 2.880 ;
        RECT  10.910 2.330 11.105 2.490 ;
        RECT  10.750 1.150 10.910 2.490 ;
        RECT  10.700 1.150 10.750 1.310 ;
        RECT  10.465 2.075 10.565 2.235 ;
        RECT  10.305 1.150 10.465 2.235 ;
        RECT  10.190 1.150 10.305 1.310 ;
        RECT  9.960 2.210 10.120 2.880 ;
        RECT  9.930 2.210 9.960 2.370 ;
        RECT  9.770 1.150 9.930 2.370 ;
        RECT  9.305 2.720 9.780 2.880 ;
        RECT  9.220 1.150 9.770 1.310 ;
        RECT  8.310 2.210 9.770 2.370 ;
        RECT  8.490 1.840 9.340 2.000 ;
        RECT  9.145 2.605 9.305 2.880 ;
        RECT  5.965 2.605 9.145 2.765 ;
        RECT  8.760 2.945 8.920 3.220 ;
        RECT  6.780 2.945 8.760 3.105 ;
        RECT  8.490 1.150 8.540 1.310 ;
        RECT  8.330 1.150 8.490 2.000 ;
        RECT  8.280 1.150 8.330 1.310 ;
        RECT  8.075 1.840 8.330 2.000 ;
        RECT  7.915 1.840 8.075 2.425 ;
        RECT  7.365 2.265 7.915 2.425 ;
        RECT  7.280 1.150 7.540 1.380 ;
        RECT  7.050 1.220 7.280 1.380 ;
        RECT  6.890 1.220 7.050 1.425 ;
        RECT  6.515 1.265 6.890 1.425 ;
        RECT  6.620 2.945 6.780 3.220 ;
        RECT  6.550 0.810 6.710 1.085 ;
        RECT  2.290 3.060 6.620 3.220 ;
        RECT  6.515 1.920 6.615 2.080 ;
        RECT  5.555 0.925 6.550 1.085 ;
        RECT  6.355 1.265 6.515 2.080 ;
        RECT  6.210 0.470 6.370 0.745 ;
        RECT  6.045 1.265 6.355 1.425 ;
        RECT  4.195 0.585 6.210 0.745 ;
        RECT  5.835 1.265 6.045 1.775 ;
        RECT  5.805 2.605 5.965 2.880 ;
        RECT  5.785 1.515 5.835 1.775 ;
        RECT  2.885 2.720 5.805 2.880 ;
        RECT  5.555 1.920 5.675 2.080 ;
        RECT  5.395 0.925 5.555 2.080 ;
        RECT  5.230 0.925 5.395 1.185 ;
        RECT  4.710 2.180 4.875 2.540 ;
        RECT  4.550 1.065 4.710 2.540 ;
        RECT  4.375 1.065 4.550 1.325 ;
        RECT  3.225 2.380 4.550 2.540 ;
        RECT  4.195 2.035 4.370 2.195 ;
        RECT  4.035 0.585 4.195 2.195 ;
        RECT  3.865 0.910 4.035 1.170 ;
        RECT  3.565 2.035 3.855 2.195 ;
        RECT  3.405 0.470 3.565 2.195 ;
        RECT  2.205 0.470 3.405 0.630 ;
        RECT  3.065 0.810 3.225 2.540 ;
        RECT  2.545 0.810 3.065 0.970 ;
        RECT  2.725 1.150 2.885 2.880 ;
        RECT  2.625 2.280 2.725 2.880 ;
        RECT  2.385 0.810 2.545 1.185 ;
        RECT  2.345 0.925 2.385 1.185 ;
        RECT  2.185 0.925 2.345 2.605 ;
        RECT  2.130 2.940 2.290 3.220 ;
        RECT  2.045 0.470 2.205 0.745 ;
        RECT  2.155 0.925 2.185 1.185 ;
        RECT  2.085 2.345 2.185 2.605 ;
        RECT  1.405 2.940 2.130 3.100 ;
        RECT  1.810 0.585 2.045 0.745 ;
        RECT  1.810 1.635 1.850 1.895 ;
        RECT  1.650 0.585 1.810 1.895 ;
        RECT  0.385 0.585 1.650 0.745 ;
        RECT  1.590 1.635 1.650 1.895 ;
        RECT  1.405 1.035 1.465 1.295 ;
        RECT  1.245 1.035 1.405 3.100 ;
        RECT  1.205 1.035 1.245 1.295 ;
        RECT  1.145 1.955 1.245 2.555 ;
        RECT  0.285 0.585 0.385 1.185 ;
        RECT  0.285 2.105 0.385 3.045 ;
        RECT  0.125 0.585 0.285 3.045 ;
    END
END AFCSHCINX4

MACRO AFCSHCINX2
    CLASS CORE ;
    FOREIGN AFCSHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.700 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.415 0.585 20.575 3.130 ;
        RECT  20.390 0.585 20.415 1.355 ;
        RECT  20.390 1.925 20.415 3.130 ;
        RECT  20.315 0.585 20.390 1.185 ;
        RECT  20.315 2.040 20.390 3.130 ;
        END
        ANTENNADIFFAREA     0.7344 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.905 0.880 20.115 1.170 ;
        RECT  19.785 1.010 19.905 1.170 ;
        RECT  19.625 1.010 19.785 1.805 ;
        RECT  19.525 1.545 19.625 1.805 ;
        END
        ANTENNAGATEAREA     0.2977 ;
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.005 0.935 13.380 1.820 ;
        RECT  12.955 1.660 13.005 1.820 ;
        RECT  12.795 1.660 12.955 2.965 ;
        END
        ANTENNADIFFAREA     0.6831 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.185 1.150 11.255 1.310 ;
        RECT  10.995 1.150 11.185 2.770 ;
        RECT  10.895 1.700 10.995 2.770 ;
        RECT  10.705 1.700 10.895 1.990 ;
        END
        ANTENNADIFFAREA     0.9460 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.465 1.700 15.975 1.990 ;
        END
        ANTENNAGATEAREA     0.4654 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.585 7.735 1.990 ;
        RECT  7.135 1.585 7.485 1.845 ;
        END
        ANTENNAGATEAREA     0.4316 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 1.290 5.595 1.645 ;
        END
        ANTENNAGATEAREA     0.7202 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.585 0.500 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.065 -0.250 20.700 0.250 ;
        RECT  19.805 -0.250 20.065 0.685 ;
        RECT  19.335 -0.250 19.805 0.250 ;
        RECT  19.175 -0.250 19.335 0.785 ;
        RECT  16.890 -0.250 19.175 0.250 ;
        RECT  15.950 -0.250 16.890 0.405 ;
        RECT  9.070 -0.250 15.950 0.250 ;
        RECT  8.810 -0.250 9.070 0.590 ;
        RECT  7.795 -0.250 8.810 0.250 ;
        RECT  7.535 -0.250 7.795 0.575 ;
        RECT  5.930 -0.250 7.535 0.250 ;
        RECT  5.670 -0.250 5.930 0.405 ;
        RECT  1.865 -0.250 5.670 0.250 ;
        RECT  1.605 -0.250 1.865 0.405 ;
        RECT  0.925 -0.250 1.605 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.065 3.440 20.700 3.940 ;
        RECT  19.805 2.955 20.065 3.940 ;
        RECT  19.245 3.440 19.805 3.940 ;
        RECT  18.985 3.115 19.245 3.940 ;
        RECT  17.005 3.440 18.985 3.940 ;
        RECT  16.745 2.260 17.005 3.940 ;
        RECT  15.445 3.440 16.745 3.940 ;
        RECT  15.185 3.285 15.445 3.940 ;
        RECT  8.535 3.440 15.185 3.940 ;
        RECT  8.275 3.100 8.535 3.940 ;
        RECT  7.545 3.440 8.275 3.940 ;
        RECT  7.285 3.100 7.545 3.940 ;
        RECT  5.945 3.440 7.285 3.940 ;
        RECT  5.685 3.285 5.945 3.940 ;
        RECT  1.915 3.440 5.685 3.940 ;
        RECT  1.655 3.285 1.915 3.940 ;
        RECT  0.895 3.440 1.655 3.940 ;
        RECT  0.635 2.595 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.135 1.585 20.215 1.845 ;
        RECT  19.975 1.585 20.135 2.680 ;
        RECT  19.335 2.520 19.975 2.680 ;
        RECT  19.335 2.170 19.615 2.330 ;
        RECT  19.335 1.035 19.445 1.295 ;
        RECT  19.175 1.035 19.335 2.330 ;
        RECT  19.175 2.520 19.335 2.935 ;
        RECT  18.995 2.170 19.175 2.330 ;
        RECT  17.975 2.775 19.175 2.935 ;
        RECT  18.835 0.585 18.995 1.805 ;
        RECT  18.835 2.170 18.995 2.595 ;
        RECT  12.275 0.585 18.835 0.745 ;
        RECT  18.315 2.435 18.835 2.595 ;
        RECT  18.495 1.035 18.655 2.255 ;
        RECT  18.275 1.035 18.495 1.295 ;
        RECT  18.155 1.555 18.315 2.595 ;
        RECT  17.975 1.035 18.025 1.295 ;
        RECT  17.815 1.035 17.975 3.200 ;
        RECT  17.765 1.035 17.815 1.295 ;
        RECT  17.465 2.260 17.515 3.200 ;
        RECT  17.305 1.035 17.465 3.200 ;
        RECT  17.255 2.260 17.305 3.200 ;
        RECT  16.965 0.925 17.125 2.005 ;
        RECT  14.395 0.925 16.965 1.085 ;
        RECT  16.445 1.265 16.495 1.425 ;
        RECT  16.445 2.385 16.495 2.985 ;
        RECT  16.285 1.265 16.445 2.985 ;
        RECT  16.235 1.265 16.285 1.425 ;
        RECT  16.235 2.385 16.285 2.985 ;
        RECT  13.515 2.780 16.235 2.940 ;
        RECT  15.725 1.265 15.985 1.520 ;
        RECT  15.275 2.205 15.985 2.365 ;
        RECT  15.275 1.360 15.725 1.520 ;
        RECT  15.115 1.360 15.275 2.365 ;
        RECT  15.035 1.745 15.115 2.005 ;
        RECT  14.805 1.265 14.935 1.425 ;
        RECT  14.805 2.270 14.855 2.530 ;
        RECT  14.645 1.265 14.805 2.530 ;
        RECT  14.235 0.925 14.395 2.600 ;
        RECT  14.135 0.925 14.235 1.250 ;
        RECT  13.780 2.340 14.235 2.600 ;
        RECT  13.785 0.935 13.885 1.195 ;
        RECT  13.625 0.935 13.785 2.160 ;
        RECT  13.515 2.000 13.625 2.160 ;
        RECT  13.355 2.000 13.515 2.940 ;
        RECT  13.255 2.270 13.355 2.940 ;
        RECT  12.655 0.975 12.815 1.235 ;
        RECT  12.615 1.075 12.655 1.235 ;
        RECT  12.455 1.075 12.615 3.135 ;
        RECT  8.875 2.975 12.455 3.135 ;
        RECT  12.115 0.585 12.275 2.770 ;
        RECT  11.525 2.610 12.115 2.770 ;
        RECT  11.890 0.470 11.935 2.035 ;
        RECT  11.775 0.470 11.890 2.430 ;
        RECT  9.845 0.470 11.775 0.630 ;
        RECT  11.730 1.875 11.775 2.430 ;
        RECT  11.525 0.810 11.595 1.695 ;
        RECT  11.435 0.810 11.525 2.770 ;
        RECT  10.185 0.810 11.435 0.970 ;
        RECT  11.365 1.535 11.435 2.770 ;
        RECT  10.525 1.150 10.745 1.310 ;
        RECT  10.525 2.170 10.675 2.795 ;
        RECT  10.365 1.150 10.525 2.795 ;
        RECT  9.220 2.635 10.365 2.795 ;
        RECT  10.025 0.810 10.185 2.450 ;
        RECT  9.865 2.190 10.025 2.450 ;
        RECT  9.685 0.470 9.845 0.930 ;
        RECT  6.615 0.770 9.685 0.930 ;
        RECT  9.515 1.155 9.675 2.455 ;
        RECT  9.405 2.195 9.515 2.455 ;
        RECT  9.175 1.765 9.335 2.025 ;
        RECT  9.060 2.415 9.220 2.795 ;
        RECT  8.335 1.815 9.175 1.975 ;
        RECT  7.160 2.415 9.060 2.575 ;
        RECT  8.715 2.755 8.875 3.135 ;
        RECT  7.095 2.755 8.715 2.915 ;
        RECT  8.175 1.115 8.335 2.235 ;
        RECT  8.075 1.115 8.175 1.275 ;
        RECT  7.945 2.075 8.175 2.235 ;
        RECT  6.955 1.115 7.255 1.275 ;
        RECT  7.000 2.065 7.160 2.575 ;
        RECT  6.935 2.755 7.095 3.105 ;
        RECT  6.955 2.065 7.000 2.325 ;
        RECT  6.795 1.115 6.955 2.325 ;
        RECT  5.495 2.945 6.935 3.105 ;
        RECT  6.275 0.430 6.885 0.590 ;
        RECT  6.745 2.065 6.795 2.325 ;
        RECT  6.485 2.505 6.745 2.765 ;
        RECT  6.495 0.770 6.615 1.275 ;
        RECT  6.455 0.770 6.495 2.255 ;
        RECT  5.155 2.605 6.485 2.765 ;
        RECT  6.335 1.015 6.455 2.255 ;
        RECT  6.255 1.015 6.335 1.275 ;
        RECT  6.235 1.995 6.335 2.255 ;
        RECT  6.115 0.430 6.275 0.745 ;
        RECT  4.275 0.585 6.115 0.745 ;
        RECT  5.935 1.495 6.085 1.755 ;
        RECT  5.775 0.925 5.935 1.985 ;
        RECT  5.130 0.925 5.775 1.085 ;
        RECT  5.405 1.825 5.775 1.985 ;
        RECT  5.335 2.945 5.495 3.220 ;
        RECT  5.145 1.825 5.405 2.255 ;
        RECT  2.260 3.060 5.335 3.220 ;
        RECT  4.995 2.605 5.155 2.875 ;
        RECT  5.005 1.825 5.145 1.985 ;
        RECT  4.845 1.475 5.005 1.985 ;
        RECT  2.965 2.715 4.995 2.875 ;
        RECT  4.665 2.190 4.815 2.535 ;
        RECT  4.665 0.960 4.715 1.220 ;
        RECT  4.505 0.960 4.665 2.535 ;
        RECT  4.455 0.960 4.505 1.220 ;
        RECT  3.305 2.375 4.505 2.535 ;
        RECT  4.275 2.035 4.325 2.195 ;
        RECT  4.115 0.585 4.275 2.195 ;
        RECT  3.945 0.585 4.115 1.305 ;
        RECT  4.065 2.035 4.115 2.195 ;
        RECT  3.645 2.035 3.815 2.195 ;
        RECT  3.485 0.470 3.645 2.195 ;
        RECT  2.205 0.470 3.485 0.630 ;
        RECT  3.145 0.810 3.305 2.535 ;
        RECT  2.545 0.810 3.145 0.970 ;
        RECT  2.885 2.195 2.965 2.875 ;
        RECT  2.725 1.150 2.885 2.875 ;
        RECT  2.705 2.195 2.725 2.875 ;
        RECT  2.455 0.810 2.545 1.240 ;
        RECT  2.385 0.810 2.455 2.595 ;
        RECT  2.295 1.030 2.385 2.595 ;
        RECT  2.165 1.030 2.295 1.290 ;
        RECT  2.195 2.335 2.295 2.595 ;
        RECT  2.100 2.940 2.260 3.220 ;
        RECT  2.045 0.470 2.205 0.785 ;
        RECT  1.970 1.665 2.115 1.925 ;
        RECT  1.405 2.940 2.100 3.100 ;
        RECT  1.970 0.625 2.045 0.785 ;
        RECT  1.810 0.625 1.970 1.925 ;
        RECT  0.385 0.625 1.810 0.785 ;
        RECT  1.405 1.035 1.465 1.295 ;
        RECT  1.145 1.035 1.405 3.100 ;
        RECT  0.680 1.245 0.840 2.330 ;
        RECT  0.385 1.245 0.680 1.405 ;
        RECT  0.385 2.170 0.680 2.330 ;
        RECT  0.125 0.585 0.385 1.405 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END AFCSHCINX2

MACRO AHHCONX4
    CLASS CORE ;
    FOREIGN AHHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.625 2.620 3.885 2.880 ;
        RECT  2.865 2.720 3.625 2.880 ;
        RECT  2.635 2.280 2.865 2.880 ;
        RECT  2.605 1.700 2.635 2.880 ;
        RECT  2.475 1.700 2.605 2.440 ;
        RECT  2.425 1.035 2.475 2.440 ;
        RECT  2.315 1.035 2.425 1.860 ;
        RECT  1.845 2.280 2.425 2.440 ;
        RECT  1.585 2.280 1.845 2.540 ;
        END
        ANTENNADIFFAREA     1.1030 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.675 0.850 6.935 2.415 ;
        RECT  4.535 0.850 6.675 1.110 ;
        RECT  6.355 2.155 6.675 2.415 ;
        RECT  6.095 2.155 6.355 3.110 ;
        RECT  5.395 2.155 6.095 2.415 ;
        RECT  5.185 2.155 5.395 3.220 ;
        RECT  5.045 2.155 5.185 3.110 ;
        END
        ANTENNADIFFAREA     1.4184 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.395 1.585 6.495 1.960 ;
        RECT  6.315 1.355 6.395 1.960 ;
        RECT  6.235 1.290 6.315 1.960 ;
        RECT  6.105 1.290 6.235 1.580 ;
        RECT  4.935 1.800 6.235 1.960 ;
        RECT  4.835 1.635 4.935 1.960 ;
        RECT  4.675 1.635 4.835 2.730 ;
        RECT  4.225 2.570 4.675 2.730 ;
        RECT  4.065 2.570 4.225 3.220 ;
        RECT  1.925 3.060 4.065 3.220 ;
        END
        ANTENNAGATEAREA     1.0075 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.545 1.455 5.645 1.615 ;
        RECT  5.370 1.290 5.545 1.615 ;
        RECT  4.290 1.290 5.370 1.450 ;
        RECT  4.145 1.290 4.290 1.590 ;
        RECT  3.885 1.290 4.145 1.825 ;
        RECT  3.805 1.290 3.885 1.580 ;
        END
        ANTENNAGATEAREA     0.8944 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.215 -0.250 7.360 0.250 ;
        RECT  6.955 -0.250 7.215 0.405 ;
        RECT  5.505 -0.250 6.955 0.250 ;
        RECT  5.245 -0.250 5.505 0.405 ;
        RECT  3.920 -0.250 5.245 0.250 ;
        RECT  3.320 -0.250 3.920 0.945 ;
        RECT  0.925 -0.250 3.320 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.875 3.440 7.360 3.940 ;
        RECT  6.615 2.595 6.875 3.940 ;
        RECT  5.845 3.440 6.615 3.940 ;
        RECT  5.585 2.595 5.845 3.940 ;
        RECT  4.795 3.440 5.585 3.940 ;
        RECT  4.535 2.935 4.795 3.940 ;
        RECT  0.925 3.440 4.535 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.025 2.110 4.285 2.370 ;
        RECT  3.375 2.210 4.025 2.370 ;
        RECT  3.275 2.210 3.375 2.540 ;
        RECT  3.115 1.195 3.275 2.540 ;
        RECT  3.035 1.195 3.115 1.355 ;
        RECT  2.775 0.695 3.035 1.355 ;
        RECT  2.135 0.695 2.775 0.855 ;
        RECT  2.095 2.620 2.355 2.880 ;
        RECT  1.975 0.695 2.135 1.430 ;
        RECT  0.385 2.720 2.095 2.880 ;
        RECT  0.985 1.270 1.975 1.430 ;
        RECT  1.335 1.625 1.830 1.785 ;
        RECT  1.635 0.585 1.795 1.030 ;
        RECT  0.285 0.585 1.635 0.745 ;
        RECT  0.625 0.925 1.335 1.085 ;
        RECT  1.175 1.625 1.335 2.515 ;
        RECT  1.075 2.255 1.175 2.515 ;
        RECT  0.625 2.255 1.075 2.415 ;
        RECT  0.825 1.270 0.985 1.825 ;
        RECT  0.465 0.925 0.625 2.415 ;
        RECT  0.285 2.595 0.385 3.195 ;
        RECT  0.125 0.585 0.285 3.195 ;
    END
END AHHCONX4

MACRO AHHCONX2
    CLASS CORE ;
    FOREIGN AHHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.625 2.620 3.885 2.880 ;
        RECT  2.865 2.720 3.625 2.880 ;
        RECT  2.640 2.280 2.865 2.880 ;
        RECT  2.605 1.770 2.640 2.880 ;
        RECT  2.475 1.770 2.605 2.440 ;
        RECT  2.315 1.035 2.475 2.440 ;
        RECT  2.140 2.110 2.315 2.440 ;
        RECT  1.845 2.280 2.140 2.440 ;
        RECT  1.585 2.280 1.845 2.540 ;
        END
        ANTENNADIFFAREA     1.1030 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.625 0.950 5.855 2.005 ;
        RECT  4.795 0.950 5.625 1.110 ;
        RECT  5.395 1.845 5.625 2.005 ;
        RECT  5.305 1.845 5.395 2.675 ;
        RECT  5.235 1.845 5.305 3.110 ;
        RECT  5.145 2.110 5.235 3.110 ;
        RECT  5.045 2.170 5.145 3.110 ;
        RECT  4.535 0.850 4.795 1.110 ;
        END
        ANTENNADIFFAREA     0.7068 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 1.635 4.935 1.990 ;
        RECT  4.675 1.635 4.835 2.730 ;
        RECT  4.225 2.570 4.675 2.730 ;
        RECT  4.065 2.570 4.225 3.220 ;
        RECT  1.925 3.060 4.065 3.220 ;
        END
        ANTENNAGATEAREA     0.7007 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.345 1.405 5.445 1.665 ;
        RECT  5.185 1.290 5.345 1.665 ;
        RECT  4.305 1.290 5.185 1.450 ;
        RECT  4.145 1.290 4.305 1.580 ;
        RECT  3.885 1.290 4.145 1.825 ;
        RECT  3.805 1.290 3.885 1.580 ;
        END
        ANTENNAGATEAREA     0.5876 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.645 -0.250 5.980 0.250 ;
        RECT  5.385 -0.250 5.645 0.750 ;
        RECT  3.925 -0.250 5.385 0.250 ;
        RECT  3.325 -0.250 3.925 1.015 ;
        RECT  0.925 -0.250 3.325 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.835 3.440 5.980 3.940 ;
        RECT  5.575 2.255 5.835 3.940 ;
        RECT  4.795 3.440 5.575 3.940 ;
        RECT  4.535 2.935 4.795 3.940 ;
        RECT  0.925 3.440 4.535 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.025 2.110 4.285 2.370 ;
        RECT  3.375 2.210 4.025 2.370 ;
        RECT  3.275 2.210 3.375 2.540 ;
        RECT  3.115 1.195 3.275 2.540 ;
        RECT  3.035 1.195 3.115 1.355 ;
        RECT  2.775 0.695 3.035 1.355 ;
        RECT  2.135 0.695 2.775 0.855 ;
        RECT  2.095 2.620 2.355 2.880 ;
        RECT  1.975 0.695 2.135 1.430 ;
        RECT  0.385 2.720 2.095 2.880 ;
        RECT  0.985 1.270 1.975 1.430 ;
        RECT  1.335 1.625 1.830 1.785 ;
        RECT  1.635 0.585 1.795 1.030 ;
        RECT  0.285 0.585 1.635 0.745 ;
        RECT  0.625 0.925 1.335 1.085 ;
        RECT  1.175 1.625 1.335 2.515 ;
        RECT  1.075 2.255 1.175 2.515 ;
        RECT  0.625 2.255 1.075 2.415 ;
        RECT  0.825 1.270 0.985 1.825 ;
        RECT  0.465 0.925 0.625 2.415 ;
        RECT  0.285 2.595 0.385 3.195 ;
        RECT  0.125 0.585 0.285 3.195 ;
    END
END AHHCONX2

MACRO AHHCINX4
    CLASS CORE ;
    FOREIGN AHHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 2.180 2.865 2.880 ;
        RECT  2.605 0.935 2.635 2.880 ;
        RECT  2.315 0.935 2.605 2.440 ;
        RECT  1.845 2.180 2.315 2.440 ;
        RECT  1.585 2.180 1.845 2.540 ;
        END
        ANTENNADIFFAREA     1.1120 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.035 7.695 3.220 ;
        RECT  7.445 1.035 7.485 3.160 ;
        RECT  6.665 1.035 7.445 1.235 ;
        RECT  7.225 2.220 7.445 3.160 ;
        RECT  5.855 2.220 7.225 2.420 ;
        RECT  6.405 0.635 6.665 1.235 ;
        RECT  5.140 0.975 6.405 1.235 ;
        RECT  5.585 2.220 5.855 3.160 ;
        RECT  4.880 0.635 5.140 1.235 ;
        END
        ANTENNADIFFAREA     1.5084 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.335 1.775 6.835 1.935 ;
        RECT  6.175 1.775 6.335 2.015 ;
        RECT  4.945 1.855 6.175 2.015 ;
        RECT  4.935 1.775 4.945 2.015 ;
        RECT  4.685 1.775 4.935 2.630 ;
        RECT  3.395 2.400 4.685 2.630 ;
        RECT  3.170 2.400 3.395 3.220 ;
        RECT  1.445 3.060 3.170 3.220 ;
        END
        ANTENNAGATEAREA     1.0504 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.585 1.465 3.865 1.625 ;
        RECT  3.265 1.275 3.585 1.625 ;
        END
        ANTENNAGATEAREA     0.5356 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.245 -0.250 7.820 0.250 ;
        RECT  6.985 -0.250 7.245 0.795 ;
        RECT  5.910 -0.250 6.985 0.250 ;
        RECT  5.910 0.535 6.080 0.795 ;
        RECT  5.650 -0.250 5.910 0.795 ;
        RECT  4.605 -0.250 5.650 0.250 ;
        RECT  5.480 0.535 5.650 0.795 ;
        RECT  4.345 -0.250 4.605 0.755 ;
        RECT  3.615 -0.250 4.345 0.250 ;
        RECT  3.355 -0.250 3.615 1.095 ;
        RECT  0.935 -0.250 3.355 0.250 ;
        RECT  0.675 -0.250 0.935 0.405 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.665 3.440 7.820 3.940 ;
        RECT  6.405 2.615 6.665 3.940 ;
        RECT  4.995 3.440 6.405 3.940 ;
        RECT  4.735 2.865 4.995 3.940 ;
        RECT  3.915 3.440 4.735 3.940 ;
        RECT  3.655 2.865 3.915 3.940 ;
        RECT  0.925 3.440 3.655 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.105 1.415 7.265 1.985 ;
        RECT  5.845 1.415 7.105 1.575 ;
        RECT  5.245 1.415 5.845 1.675 ;
        RECT  4.465 1.415 5.245 1.575 ;
        RECT  4.205 1.005 4.465 2.215 ;
        RECT  3.905 1.005 4.205 1.265 ;
        RECT  3.115 1.840 3.375 2.215 ;
        RECT  3.085 1.840 3.115 2.000 ;
        RECT  2.925 0.595 3.085 2.000 ;
        RECT  2.825 0.595 2.925 1.195 ;
        RECT  2.135 0.595 2.825 0.755 ;
        RECT  2.095 2.620 2.355 2.880 ;
        RECT  1.975 0.595 2.135 1.545 ;
        RECT  1.875 1.740 2.135 2.000 ;
        RECT  0.385 2.720 2.095 2.880 ;
        RECT  0.965 1.385 1.975 1.545 ;
        RECT  1.335 1.840 1.875 2.000 ;
        RECT  1.635 0.585 1.795 1.190 ;
        RECT  0.285 0.585 1.635 0.745 ;
        RECT  0.625 0.925 1.335 1.085 ;
        RECT  1.175 1.840 1.335 2.520 ;
        RECT  1.075 2.095 1.175 2.520 ;
        RECT  0.625 2.095 1.075 2.255 ;
        RECT  0.805 1.385 0.965 1.825 ;
        RECT  0.465 0.925 0.625 2.255 ;
        RECT  0.285 2.595 0.385 3.195 ;
        RECT  0.125 0.585 0.285 3.195 ;
    END
END AHHCINX4

MACRO AHHCINX2
    CLASS CORE ;
    FOREIGN AHHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 2.280 2.865 2.880 ;
        RECT  2.605 1.035 2.635 2.880 ;
        RECT  2.415 1.035 2.605 2.440 ;
        RECT  2.315 1.035 2.415 1.295 ;
        RECT  1.845 2.280 2.415 2.440 ;
        RECT  1.585 2.280 1.845 2.540 ;
        END
        ANTENNADIFFAREA     1.1120 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.375 2.095 4.635 2.695 ;
        RECT  4.365 2.095 4.375 2.400 ;
        RECT  4.265 1.065 4.365 2.400 ;
        RECT  4.205 1.065 4.265 2.255 ;
        RECT  4.195 1.065 4.205 1.225 ;
        RECT  3.935 0.965 4.195 1.225 ;
        END
        ANTENNADIFFAREA     0.6572 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.075 1.585 5.235 3.035 ;
        RECT  4.015 2.875 5.075 3.035 ;
        RECT  4.015 1.405 4.025 1.665 ;
        RECT  3.805 1.405 4.015 3.035 ;
        RECT  3.765 1.405 3.805 1.665 ;
        RECT  3.370 2.875 3.805 3.035 ;
        RECT  3.200 2.875 3.370 3.220 ;
        RECT  1.445 3.060 3.200 3.220 ;
        END
        ANTENNAGATEAREA     0.7163 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.210 0.475 5.455 0.635 ;
        RECT  5.035 0.475 5.210 0.745 ;
        RECT  3.555 0.585 5.035 0.745 ;
        RECT  3.530 1.170 3.560 1.755 ;
        RECT  3.530 0.585 3.555 0.880 ;
        RECT  3.370 0.585 3.530 1.755 ;
        RECT  3.345 1.170 3.370 1.755 ;
        RECT  3.285 1.290 3.345 1.755 ;
        END
        ANTENNAGATEAREA     0.4056 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.735 -0.250 5.980 0.250 ;
        RECT  4.475 -0.250 4.735 0.405 ;
        RECT  3.640 -0.250 4.475 0.250 ;
        RECT  3.380 -0.250 3.640 0.405 ;
        RECT  0.925 -0.250 3.380 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.345 3.440 5.980 3.940 ;
        RECT  5.085 3.285 5.345 3.940 ;
        RECT  3.925 3.440 5.085 3.940 ;
        RECT  3.665 3.285 3.925 3.940 ;
        RECT  0.925 3.440 3.665 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.595 2.835 5.855 3.095 ;
        RECT  5.575 2.835 5.595 2.995 ;
        RECT  5.415 0.895 5.575 2.995 ;
        RECT  4.805 1.245 5.415 1.405 ;
        RECT  4.645 1.245 4.805 1.675 ;
        RECT  4.545 1.415 4.645 1.675 ;
        RECT  3.115 1.940 3.375 2.555 ;
        RECT  3.085 1.940 3.115 2.100 ;
        RECT  2.925 0.585 3.085 2.100 ;
        RECT  2.825 0.585 2.925 1.185 ;
        RECT  2.135 0.585 2.825 0.745 ;
        RECT  2.095 2.620 2.355 2.880 ;
        RECT  1.975 0.585 2.135 1.640 ;
        RECT  1.875 1.830 2.135 2.090 ;
        RECT  0.385 2.720 2.095 2.880 ;
        RECT  0.985 1.480 1.975 1.640 ;
        RECT  1.335 1.930 1.875 2.090 ;
        RECT  1.635 0.585 1.795 1.185 ;
        RECT  0.285 0.585 1.635 0.745 ;
        RECT  0.625 0.925 1.335 1.085 ;
        RECT  1.175 1.930 1.335 2.515 ;
        RECT  1.075 2.255 1.175 2.515 ;
        RECT  0.625 2.255 1.075 2.415 ;
        RECT  0.825 1.480 0.985 1.825 ;
        RECT  0.465 0.925 0.625 2.415 ;
        RECT  0.285 2.595 0.385 3.195 ;
        RECT  0.125 0.585 0.285 3.195 ;
    END
END AHHCINX2

MACRO ACHCONX4
    CLASS CORE ;
    FOREIGN ACHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.155 0.955 8.255 1.215 ;
        RECT  7.995 0.955 8.155 2.400 ;
        RECT  7.945 1.015 7.995 2.400 ;
        RECT  7.235 1.015 7.945 1.175 ;
        RECT  7.845 2.145 7.945 2.400 ;
        RECT  7.585 2.145 7.845 2.745 ;
        RECT  6.945 2.585 7.585 2.745 ;
        RECT  6.975 0.565 7.235 1.175 ;
        RECT  6.785 2.585 6.945 3.120 ;
        RECT  6.515 2.860 6.785 3.120 ;
        END
        ANTENNADIFFAREA     1.4431 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.510 1.700 9.535 1.990 ;
        RECT  9.475 1.640 9.510 1.990 ;
        RECT  9.325 1.590 9.475 1.990 ;
        RECT  8.875 1.590 9.325 1.850 ;
        END
        ANTENNAGATEAREA     0.5226 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.645 1.290 5.855 1.775 ;
        RECT  5.255 1.515 5.645 1.775 ;
        END
        ANTENNAGATEAREA     1.0673 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.605 0.555 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 -0.250 10.120 0.250 ;
        RECT  9.585 -0.250 9.845 1.175 ;
        RECT  8.765 -0.250 9.585 0.250 ;
        RECT  8.505 -0.250 8.765 0.405 ;
        RECT  5.805 -0.250 8.505 0.250 ;
        RECT  5.545 -0.250 5.805 0.405 ;
        RECT  0.925 -0.250 5.545 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.810 3.440 10.120 3.940 ;
        RECT  9.210 2.170 9.810 3.940 ;
        RECT  8.365 3.440 9.210 3.940 ;
        RECT  8.105 3.285 8.365 3.940 ;
        RECT  5.755 3.440 8.105 3.940 ;
        RECT  5.495 2.950 5.755 3.940 ;
        RECT  0.985 3.440 5.495 3.940 ;
        RECT  0.725 2.615 0.985 3.940 ;
        RECT  0.000 3.440 0.725 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.045 0.610 9.305 1.210 ;
        RECT  8.595 0.610 9.045 0.770 ;
        RECT  8.645 2.160 8.905 3.100 ;
        RECT  8.595 2.160 8.645 2.320 ;
        RECT  7.285 2.925 8.645 3.085 ;
        RECT  8.435 0.610 8.595 2.320 ;
        RECT  7.745 0.610 8.435 0.770 ;
        RECT  7.485 0.510 7.745 0.770 ;
        RECT  7.315 1.410 7.575 1.670 ;
        RECT  6.795 1.410 7.315 1.570 ;
        RECT  7.125 2.925 7.285 3.185 ;
        RECT  6.965 1.765 7.065 2.025 ;
        RECT  6.805 1.765 6.965 2.365 ;
        RECT  6.605 2.205 6.805 2.365 ;
        RECT  6.635 0.630 6.795 1.570 ;
        RECT  4.635 0.630 6.635 0.790 ;
        RECT  6.535 1.410 6.635 1.570 ;
        RECT  6.445 2.205 6.605 2.680 ;
        RECT  6.375 1.410 6.535 1.865 ;
        RECT  6.195 0.970 6.445 1.230 ;
        RECT  5.125 2.520 6.445 2.680 ;
        RECT  6.195 2.075 6.265 2.335 ;
        RECT  6.035 0.970 6.195 2.335 ;
        RECT  6.005 2.075 6.035 2.335 ;
        RECT  5.075 2.075 5.245 2.335 ;
        RECT  5.075 1.055 5.145 1.315 ;
        RECT  4.965 2.520 5.125 3.165 ;
        RECT  4.915 1.055 5.075 2.335 ;
        RECT  1.325 3.005 4.965 3.165 ;
        RECT  4.885 1.055 4.915 1.315 ;
        RECT  4.735 1.555 4.915 1.815 ;
        RECT  4.555 2.085 4.735 2.685 ;
        RECT  4.375 0.630 4.635 1.255 ;
        RECT  4.395 1.475 4.555 2.825 ;
        RECT  4.125 1.475 4.395 1.635 ;
        RECT  1.665 2.665 4.395 2.825 ;
        RECT  3.615 0.630 4.375 0.790 ;
        RECT  4.115 2.170 4.215 2.430 ;
        RECT  3.965 0.970 4.125 1.635 ;
        RECT  3.955 1.825 4.115 2.430 ;
        RECT  3.865 0.970 3.965 1.230 ;
        RECT  3.615 1.825 3.955 1.985 ;
        RECT  3.445 2.225 3.705 2.485 ;
        RECT  3.455 0.630 3.615 1.985 ;
        RECT  3.355 0.995 3.455 1.255 ;
        RECT  2.915 2.325 3.445 2.485 ;
        RECT  2.915 0.720 3.105 1.320 ;
        RECT  2.755 0.435 2.915 2.485 ;
        RECT  2.135 0.435 2.755 0.595 ;
        RECT  2.505 2.325 2.755 2.485 ;
        RECT  2.315 0.775 2.575 1.375 ;
        RECT  1.605 0.820 2.315 0.980 ;
        RECT  1.975 0.435 2.135 0.630 ;
        RECT  1.945 1.165 2.065 1.325 ;
        RECT  1.265 0.470 1.975 0.630 ;
        RECT  1.785 1.165 1.945 2.040 ;
        RECT  1.665 1.880 1.785 2.040 ;
        RECT  1.505 1.880 1.665 2.825 ;
        RECT  1.445 0.820 1.605 1.085 ;
        RECT  1.325 0.925 1.445 1.085 ;
        RECT  1.165 0.925 1.325 3.165 ;
        RECT  1.105 0.470 1.265 0.745 ;
        RECT  0.385 0.585 1.105 0.745 ;
        RECT  0.825 1.035 0.985 2.330 ;
        RECT  0.385 1.035 0.825 1.195 ;
        RECT  0.385 2.170 0.825 2.330 ;
        RECT  0.125 0.585 0.385 1.195 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END ACHCONX4

MACRO ACHCONX2
    CLASS CORE ;
    FOREIGN ACHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.965 1.010 7.125 1.995 ;
        RECT  6.485 1.010 6.965 1.170 ;
        RECT  6.645 1.835 6.965 1.995 ;
        RECT  6.485 1.835 6.645 2.730 ;
        RECT  6.225 0.565 6.485 1.170 ;
        RECT  6.165 2.570 6.485 2.730 ;
        RECT  6.005 2.570 6.165 3.120 ;
        RECT  5.855 2.860 6.005 3.120 ;
        RECT  5.645 2.860 5.855 3.220 ;
        END
        ANTENNADIFFAREA     0.8101 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.565 2.520 7.695 2.845 ;
        RECT  7.305 2.515 7.565 2.845 ;
        END
        ANTENNAGATEAREA     0.2613 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 1.515 5.080 1.775 ;
        RECT  4.725 1.515 4.935 1.990 ;
        RECT  4.480 1.515 4.725 1.775 ;
        END
        ANTENNAGATEAREA     0.9854 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.605 0.555 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.605 -0.250 7.820 0.250 ;
        RECT  7.345 -0.250 7.605 0.405 ;
        RECT  5.135 -0.250 7.345 0.250 ;
        RECT  4.875 -0.250 5.135 0.405 ;
        RECT  0.925 -0.250 4.875 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.205 3.440 7.820 3.940 ;
        RECT  6.945 3.285 7.205 3.940 ;
        RECT  4.940 3.440 6.945 3.940 ;
        RECT  4.680 2.950 4.940 3.940 ;
        RECT  0.985 3.440 4.680 3.940 ;
        RECT  0.725 2.615 0.985 3.940 ;
        RECT  0.000 3.440 0.725 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.305 0.660 7.465 2.335 ;
        RECT  7.005 0.660 7.305 0.820 ;
        RECT  7.000 2.175 7.305 2.335 ;
        RECT  6.745 0.560 7.005 0.820 ;
        RECT  6.840 2.175 7.000 3.075 ;
        RECT  6.605 2.915 6.840 3.075 ;
        RECT  6.625 1.350 6.785 1.645 ;
        RECT  5.965 1.350 6.625 1.510 ;
        RECT  6.345 2.915 6.605 3.175 ;
        RECT  6.145 1.690 6.305 2.365 ;
        RECT  5.825 2.205 6.145 2.365 ;
        RECT  5.805 0.640 5.965 1.865 ;
        RECT  5.665 2.205 5.825 2.680 ;
        RECT  4.485 0.640 5.805 0.800 ;
        RECT  5.610 1.605 5.805 1.865 ;
        RECT  4.205 2.520 5.665 2.680 ;
        RECT  5.465 1.025 5.625 1.350 ;
        RECT  5.430 2.075 5.480 2.335 ;
        RECT  5.430 1.190 5.465 1.350 ;
        RECT  5.270 1.190 5.430 2.335 ;
        RECT  5.220 2.075 5.270 2.335 ;
        RECT  4.335 1.055 4.595 1.330 ;
        RECT  4.325 0.470 4.485 0.800 ;
        RECT  4.205 2.075 4.400 2.335 ;
        RECT  4.205 1.170 4.335 1.330 ;
        RECT  3.525 0.470 4.325 0.630 ;
        RECT  4.045 1.170 4.205 2.335 ;
        RECT  4.045 2.520 4.205 3.185 ;
        RECT  3.865 0.810 4.085 0.970 ;
        RECT  1.325 3.025 4.045 3.185 ;
        RECT  3.705 0.810 3.865 2.845 ;
        RECT  3.555 2.585 3.705 2.845 ;
        RECT  1.665 2.685 3.555 2.845 ;
        RECT  3.365 0.470 3.525 2.405 ;
        RECT  3.305 2.245 3.365 2.405 ;
        RECT  3.045 2.245 3.305 2.505 ;
        RECT  2.965 0.685 3.065 1.285 ;
        RECT  2.805 0.470 2.965 1.880 ;
        RECT  1.265 0.470 2.805 0.630 ;
        RECT  2.795 1.720 2.805 1.880 ;
        RECT  2.635 1.720 2.795 2.505 ;
        RECT  2.535 2.245 2.635 2.505 ;
        RECT  2.455 0.935 2.555 1.195 ;
        RECT  2.295 0.820 2.455 1.195 ;
        RECT  1.605 0.820 2.295 0.980 ;
        RECT  1.945 1.165 2.045 1.325 ;
        RECT  1.785 1.165 1.945 2.040 ;
        RECT  1.665 1.880 1.785 2.040 ;
        RECT  1.505 1.880 1.665 2.845 ;
        RECT  1.445 0.820 1.605 1.085 ;
        RECT  1.325 0.925 1.445 1.085 ;
        RECT  1.165 0.925 1.325 3.185 ;
        RECT  1.105 0.470 1.265 0.745 ;
        RECT  0.385 0.585 1.105 0.745 ;
        RECT  0.825 1.035 0.985 2.330 ;
        RECT  0.385 1.035 0.825 1.195 ;
        RECT  0.385 2.170 0.825 2.330 ;
        RECT  0.125 0.585 0.385 1.195 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END ACHCONX2

MACRO ACHCINX4
    CLASS CORE ;
    FOREIGN ACHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.155 0.955 8.315 1.215 ;
        RECT  8.055 0.955 8.155 2.400 ;
        RECT  7.945 1.015 8.055 2.400 ;
        RECT  7.295 1.015 7.945 1.175 ;
        RECT  7.845 2.145 7.945 2.400 ;
        RECT  7.585 2.145 7.845 2.745 ;
        RECT  6.945 2.585 7.585 2.745 ;
        RECT  7.025 0.565 7.295 1.175 ;
        RECT  6.785 2.585 6.945 3.120 ;
        RECT  6.515 2.860 6.785 3.120 ;
        END
        ANTENNADIFFAREA     1.4542 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.510 1.700 9.535 1.990 ;
        RECT  9.475 1.640 9.510 1.990 ;
        RECT  9.325 1.590 9.475 1.990 ;
        RECT  8.875 1.590 9.325 1.850 ;
        END
        ANTENNAGATEAREA     0.5226 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.645 2.110 5.855 2.400 ;
        RECT  5.570 2.110 5.645 2.270 ;
        RECT  5.410 1.515 5.570 2.270 ;
        RECT  5.275 1.515 5.410 1.775 ;
        END
        ANTENNAGATEAREA     0.7917 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.605 0.555 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.905 -0.250 10.120 0.250 ;
        RECT  9.645 -0.250 9.905 1.175 ;
        RECT  8.825 -0.250 9.645 0.250 ;
        RECT  8.565 -0.250 8.825 0.405 ;
        RECT  5.810 -0.250 8.565 0.250 ;
        RECT  5.550 -0.250 5.810 0.405 ;
        RECT  0.925 -0.250 5.550 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.810 3.440 10.120 3.940 ;
        RECT  9.210 2.170 9.810 3.940 ;
        RECT  8.365 3.440 9.210 3.940 ;
        RECT  8.105 3.285 8.365 3.940 ;
        RECT  5.755 3.440 8.105 3.940 ;
        RECT  5.495 2.950 5.755 3.940 ;
        RECT  0.985 3.440 5.495 3.940 ;
        RECT  0.725 2.615 0.985 3.940 ;
        RECT  0.000 3.440 0.725 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.105 0.610 9.365 1.210 ;
        RECT  8.655 0.610 9.105 0.770 ;
        RECT  8.655 2.160 8.905 3.100 ;
        RECT  8.645 0.610 8.655 3.100 ;
        RECT  8.495 0.610 8.645 2.320 ;
        RECT  7.285 2.925 8.645 3.085 ;
        RECT  7.805 0.610 8.495 0.770 ;
        RECT  7.545 0.510 7.805 0.770 ;
        RECT  7.375 1.410 7.635 1.670 ;
        RECT  6.820 1.410 7.375 1.570 ;
        RECT  7.125 2.925 7.285 3.185 ;
        RECT  7.025 1.765 7.125 2.025 ;
        RECT  6.865 1.765 7.025 2.365 ;
        RECT  6.605 2.205 6.865 2.365 ;
        RECT  6.660 0.610 6.820 1.570 ;
        RECT  4.635 0.610 6.660 0.770 ;
        RECT  6.595 1.410 6.660 1.570 ;
        RECT  6.445 2.205 6.605 2.680 ;
        RECT  6.435 1.410 6.595 1.865 ;
        RECT  6.255 0.970 6.465 1.230 ;
        RECT  6.230 2.520 6.445 2.680 ;
        RECT  6.215 0.970 6.255 2.025 ;
        RECT  6.070 2.520 6.230 2.750 ;
        RECT  6.095 0.970 6.215 2.335 ;
        RECT  6.055 1.865 6.095 2.335 ;
        RECT  5.125 2.590 6.070 2.750 ;
        RECT  5.755 1.055 5.915 1.685 ;
        RECT  5.145 1.055 5.755 1.215 ;
        RECT  5.075 2.075 5.195 2.335 ;
        RECT  5.075 1.055 5.145 1.315 ;
        RECT  4.965 2.590 5.125 3.165 ;
        RECT  4.915 1.055 5.075 2.335 ;
        RECT  1.325 3.005 4.965 3.165 ;
        RECT  4.885 1.055 4.915 1.315 ;
        RECT  4.735 1.555 4.915 1.815 ;
        RECT  4.555 2.085 4.735 2.685 ;
        RECT  4.475 0.610 4.635 1.255 ;
        RECT  4.395 1.475 4.555 2.825 ;
        RECT  4.375 0.630 4.475 1.255 ;
        RECT  4.125 1.475 4.395 1.635 ;
        RECT  1.665 2.665 4.395 2.825 ;
        RECT  3.615 0.630 4.375 0.790 ;
        RECT  4.115 2.170 4.215 2.430 ;
        RECT  3.965 0.970 4.125 1.635 ;
        RECT  3.955 1.825 4.115 2.430 ;
        RECT  3.865 0.970 3.965 1.230 ;
        RECT  3.615 1.825 3.955 1.985 ;
        RECT  3.445 2.225 3.705 2.485 ;
        RECT  3.455 0.630 3.615 1.985 ;
        RECT  3.355 0.995 3.455 1.255 ;
        RECT  2.915 2.325 3.445 2.485 ;
        RECT  2.915 0.720 3.105 1.320 ;
        RECT  2.755 0.435 2.915 2.485 ;
        RECT  2.135 0.435 2.755 0.595 ;
        RECT  2.505 2.325 2.755 2.485 ;
        RECT  2.315 0.775 2.575 1.375 ;
        RECT  1.605 0.820 2.315 0.980 ;
        RECT  1.975 0.435 2.135 0.630 ;
        RECT  1.945 1.165 2.065 1.325 ;
        RECT  1.265 0.470 1.975 0.630 ;
        RECT  1.785 1.165 1.945 2.040 ;
        RECT  1.665 1.880 1.785 2.040 ;
        RECT  1.505 1.880 1.665 2.825 ;
        RECT  1.445 0.820 1.605 1.085 ;
        RECT  1.325 0.925 1.445 1.085 ;
        RECT  1.165 0.925 1.325 3.165 ;
        RECT  1.105 0.470 1.265 0.745 ;
        RECT  0.385 0.585 1.105 0.745 ;
        RECT  0.825 1.035 0.985 2.330 ;
        RECT  0.385 1.035 0.825 1.195 ;
        RECT  0.385 2.170 0.825 2.330 ;
        RECT  0.125 0.585 0.385 1.195 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END ACHCINX4

MACRO ACHCINX2
    CLASS CORE ;
    FOREIGN ACHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.015 1.010 7.175 1.995 ;
        RECT  6.590 1.010 7.015 1.170 ;
        RECT  6.700 1.835 7.015 1.995 ;
        RECT  6.540 1.835 6.700 2.730 ;
        RECT  6.330 0.565 6.590 1.170 ;
        RECT  6.165 2.570 6.540 2.730 ;
        RECT  6.005 2.570 6.165 3.120 ;
        RECT  5.855 2.860 6.005 3.120 ;
        RECT  5.645 2.860 5.855 3.220 ;
        END
        ANTENNADIFFAREA     0.8978 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.565 2.520 7.695 2.845 ;
        RECT  7.305 2.515 7.565 2.845 ;
        END
        ANTENNAGATEAREA     0.2613 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.785 2.110 4.935 2.400 ;
        RECT  4.625 1.515 4.785 2.400 ;
        RECT  4.480 1.515 4.625 1.775 ;
        END
        ANTENNAGATEAREA     0.7098 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.605 0.555 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.695 -0.250 7.820 0.250 ;
        RECT  7.435 -0.250 7.695 0.405 ;
        RECT  5.135 -0.250 7.435 0.250 ;
        RECT  4.875 -0.250 5.135 0.405 ;
        RECT  0.925 -0.250 4.875 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.205 3.440 7.820 3.940 ;
        RECT  6.945 3.285 7.205 3.940 ;
        RECT  4.940 3.440 6.945 3.940 ;
        RECT  4.680 2.950 4.940 3.940 ;
        RECT  0.985 3.440 4.680 3.940 ;
        RECT  0.725 2.615 0.985 3.940 ;
        RECT  0.000 3.440 0.725 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.355 0.660 7.515 2.335 ;
        RECT  7.110 0.660 7.355 0.820 ;
        RECT  7.045 2.175 7.355 2.335 ;
        RECT  6.850 0.560 7.110 0.820 ;
        RECT  6.885 2.175 7.045 3.075 ;
        RECT  6.605 2.915 6.885 3.075 ;
        RECT  6.675 1.350 6.835 1.645 ;
        RECT  5.965 1.350 6.675 1.510 ;
        RECT  6.345 2.915 6.605 3.175 ;
        RECT  6.195 1.690 6.355 2.365 ;
        RECT  5.825 2.205 6.195 2.365 ;
        RECT  5.875 0.640 5.965 1.765 ;
        RECT  5.805 0.640 5.875 1.865 ;
        RECT  5.665 2.205 5.825 2.680 ;
        RECT  4.485 0.640 5.805 0.800 ;
        RECT  5.715 1.605 5.805 1.865 ;
        RECT  5.325 2.520 5.665 2.680 ;
        RECT  5.535 1.025 5.625 1.350 ;
        RECT  5.480 1.025 5.535 2.025 ;
        RECT  5.465 1.025 5.480 2.335 ;
        RECT  5.375 1.190 5.465 2.335 ;
        RECT  5.320 1.865 5.375 2.335 ;
        RECT  5.165 2.520 5.325 2.755 ;
        RECT  5.220 2.075 5.320 2.335 ;
        RECT  5.035 1.155 5.195 1.685 ;
        RECT  4.205 2.595 5.165 2.755 ;
        RECT  4.595 1.155 5.035 1.315 ;
        RECT  4.335 1.055 4.595 1.315 ;
        RECT  4.325 0.470 4.485 0.800 ;
        RECT  4.205 2.075 4.400 2.335 ;
        RECT  4.205 1.155 4.335 1.315 ;
        RECT  3.525 0.470 4.325 0.630 ;
        RECT  4.140 1.155 4.205 2.335 ;
        RECT  4.045 2.595 4.205 3.185 ;
        RECT  4.045 1.155 4.140 2.285 ;
        RECT  3.865 0.810 4.085 0.970 ;
        RECT  1.325 3.025 4.045 3.185 ;
        RECT  3.705 0.810 3.865 2.845 ;
        RECT  3.555 2.585 3.705 2.845 ;
        RECT  1.665 2.685 3.555 2.845 ;
        RECT  3.365 0.470 3.525 2.405 ;
        RECT  3.305 2.245 3.365 2.405 ;
        RECT  3.045 2.245 3.305 2.505 ;
        RECT  2.965 0.685 3.065 1.285 ;
        RECT  2.805 0.470 2.965 1.880 ;
        RECT  1.265 0.470 2.805 0.630 ;
        RECT  2.795 1.720 2.805 1.880 ;
        RECT  2.635 1.720 2.795 2.505 ;
        RECT  2.535 2.245 2.635 2.505 ;
        RECT  2.455 0.935 2.555 1.195 ;
        RECT  2.295 0.820 2.455 1.195 ;
        RECT  1.605 0.820 2.295 0.980 ;
        RECT  1.945 1.165 2.045 1.325 ;
        RECT  1.785 1.165 1.945 2.040 ;
        RECT  1.665 1.880 1.785 2.040 ;
        RECT  1.505 1.880 1.665 2.845 ;
        RECT  1.445 0.820 1.605 1.085 ;
        RECT  1.325 0.925 1.445 1.085 ;
        RECT  1.165 0.925 1.325 3.185 ;
        RECT  1.105 0.470 1.265 0.745 ;
        RECT  0.385 0.585 1.105 0.745 ;
        RECT  0.825 1.035 0.985 2.330 ;
        RECT  0.385 1.035 0.825 1.195 ;
        RECT  0.385 2.170 0.825 2.330 ;
        RECT  0.125 0.585 0.385 1.195 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END ACHCINX2

MACRO AFHCONX4
    CLASS CORE ;
    FOREIGN AFHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.800 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.515 0.655 13.675 3.055 ;
        RECT  13.415 0.655 13.515 1.255 ;
        RECT  13.465 2.110 13.515 3.055 ;
        RECT  13.415 2.115 13.465 3.055 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 0.830 7.725 0.990 ;
        RECT  6.625 2.605 7.695 2.765 ;
        RECT  6.625 0.830 6.775 1.765 ;
        RECT  6.565 0.830 6.625 2.765 ;
        RECT  6.465 0.940 6.565 2.765 ;
        RECT  6.345 0.940 6.465 1.200 ;
        END
        ANTENNADIFFAREA     1.5167 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.865 1.530 9.075 1.990 ;
        RECT  8.425 1.530 8.865 1.790 ;
        END
        ANTENNAGATEAREA     1.1024 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 1.440 5.485 1.805 ;
        RECT  5.185 1.290 5.395 1.805 ;
        RECT  5.170 1.440 5.185 1.805 ;
        END
        ANTENNAGATEAREA     1.0751 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.540 0.530 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.045 -0.250 13.800 0.250 ;
        RECT  12.785 -0.250 13.045 0.405 ;
        RECT  10.795 -0.250 12.785 0.250 ;
        RECT  10.535 -0.250 10.795 0.405 ;
        RECT  9.715 -0.250 10.535 0.250 ;
        RECT  9.455 -0.250 9.715 0.405 ;
        RECT  8.635 -0.250 9.455 0.250 ;
        RECT  8.375 -0.250 8.635 0.405 ;
        RECT  5.285 -0.250 8.375 0.250 ;
        RECT  5.025 -0.250 5.285 0.405 ;
        RECT  0.925 -0.250 5.025 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.115 3.440 13.800 3.940 ;
        RECT  12.855 3.285 13.115 3.940 ;
        RECT  10.625 3.440 12.855 3.940 ;
        RECT  10.365 3.285 10.625 3.940 ;
        RECT  9.515 3.440 10.365 3.940 ;
        RECT  9.255 3.285 9.515 3.940 ;
        RECT  8.435 3.440 9.255 3.940 ;
        RECT  8.175 3.285 8.435 3.940 ;
        RECT  5.605 3.440 8.175 3.940 ;
        RECT  5.345 3.285 5.605 3.940 ;
        RECT  1.110 3.440 5.345 3.940 ;
        RECT  0.850 2.610 1.110 3.940 ;
        RECT  0.000 3.440 0.850 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.230 1.510 13.335 1.770 ;
        RECT  13.070 1.510 13.230 3.105 ;
        RECT  12.015 2.945 13.070 3.105 ;
        RECT  12.655 0.625 12.815 1.675 ;
        RECT  12.610 0.625 12.655 0.785 ;
        RECT  12.450 0.490 12.610 0.785 ;
        RECT  12.475 2.110 12.575 2.710 ;
        RECT  12.315 0.965 12.475 2.710 ;
        RECT  11.210 0.490 12.450 0.650 ;
        RECT  12.280 0.965 12.315 1.125 ;
        RECT  12.020 0.915 12.280 1.125 ;
        RECT  12.015 1.305 12.135 2.245 ;
        RECT  11.975 1.305 12.015 3.105 ;
        RECT  11.720 1.305 11.975 1.465 ;
        RECT  11.855 2.085 11.975 3.105 ;
        RECT  11.675 1.645 11.795 1.905 ;
        RECT  11.560 0.865 11.720 1.465 ;
        RECT  11.515 1.645 11.675 3.105 ;
        RECT  8.040 2.945 11.515 3.105 ;
        RECT  11.050 0.490 11.210 2.675 ;
        RECT  10.935 2.075 11.050 2.675 ;
        RECT  10.055 2.075 10.935 2.235 ;
        RECT  10.700 0.590 10.860 1.825 ;
        RECT  8.075 0.590 10.700 0.750 ;
        RECT  10.055 0.940 10.255 1.200 ;
        RECT  9.795 0.940 10.055 2.765 ;
        RECT  9.285 1.185 9.445 2.330 ;
        RECT  9.175 1.185 9.285 1.345 ;
        RECT  8.975 2.170 9.285 2.330 ;
        RECT  8.915 0.940 9.175 1.345 ;
        RECT  8.715 2.170 8.975 2.765 ;
        RECT  8.235 1.185 8.915 1.345 ;
        RECT  7.975 0.940 8.235 1.345 ;
        RECT  7.915 0.470 8.075 0.750 ;
        RECT  7.880 1.895 8.040 3.105 ;
        RECT  7.115 1.185 7.975 1.345 ;
        RECT  6.165 0.470 7.915 0.630 ;
        RECT  7.695 1.895 7.880 2.055 ;
        RECT  4.950 2.945 7.880 3.105 ;
        RECT  7.115 2.260 7.185 2.420 ;
        RECT  6.955 1.185 7.115 2.420 ;
        RECT  6.925 2.260 6.955 2.420 ;
        RECT  6.165 1.705 6.285 1.965 ;
        RECT  6.005 0.470 6.165 1.965 ;
        RECT  5.935 2.165 6.095 2.765 ;
        RECT  4.845 0.585 6.005 0.745 ;
        RECT  5.825 2.165 5.935 2.325 ;
        RECT  5.665 0.940 5.825 2.325 ;
        RECT  5.565 0.940 5.665 1.200 ;
        RECT  4.965 2.160 5.065 2.760 ;
        RECT  4.805 1.305 4.965 2.760 ;
        RECT  4.790 2.945 4.950 3.165 ;
        RECT  4.685 0.500 4.845 0.745 ;
        RECT  4.745 1.305 4.805 1.465 ;
        RECT  2.195 3.005 4.790 3.165 ;
        RECT  4.485 0.960 4.745 1.465 ;
        RECT  4.095 0.500 4.685 0.660 ;
        RECT  4.455 2.225 4.555 2.825 ;
        RECT  3.935 1.305 4.485 1.465 ;
        RECT  4.295 1.645 4.455 2.825 ;
        RECT  3.755 1.645 4.295 1.805 ;
        RECT  2.540 2.665 4.295 2.825 ;
        RECT  3.935 0.470 4.095 0.660 ;
        RECT  3.945 2.180 4.045 2.440 ;
        RECT  3.785 1.985 3.945 2.440 ;
        RECT  3.415 0.470 3.935 0.630 ;
        RECT  3.415 1.985 3.785 2.145 ;
        RECT  3.595 0.810 3.755 1.805 ;
        RECT  3.075 2.325 3.535 2.485 ;
        RECT  3.255 0.470 3.415 2.145 ;
        RECT  3.035 0.750 3.255 1.010 ;
        RECT  2.915 1.340 3.075 2.485 ;
        RECT  2.735 1.340 2.915 1.500 ;
        RECT  2.720 2.325 2.915 2.485 ;
        RECT  2.575 0.495 2.735 1.500 ;
        RECT  1.265 0.495 2.575 0.655 ;
        RECT  2.395 1.685 2.540 2.825 ;
        RECT  2.380 0.835 2.395 2.825 ;
        RECT  2.235 0.835 2.380 1.845 ;
        RECT  1.605 0.835 2.235 0.995 ;
        RECT  2.055 2.335 2.195 3.165 ;
        RECT  2.030 1.175 2.055 3.165 ;
        RECT  1.895 1.175 2.030 2.935 ;
        RECT  1.605 2.175 1.685 3.115 ;
        RECT  1.445 0.835 1.605 3.115 ;
        RECT  1.305 1.025 1.445 1.285 ;
        RECT  1.425 2.175 1.445 3.115 ;
        RECT  1.105 0.495 1.265 0.755 ;
        RECT  1.015 1.470 1.215 1.730 ;
        RECT  0.385 0.595 1.105 0.755 ;
        RECT  0.855 1.035 1.015 2.330 ;
        RECT  0.385 1.035 0.855 1.195 ;
        RECT  0.560 2.170 0.855 2.330 ;
        RECT  0.300 2.170 0.560 3.110 ;
        RECT  0.125 0.595 0.385 1.195 ;
    END
END AFHCONX4

MACRO AFHCONX2
    CLASS CORE ;
    FOREIGN AFHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.165 0.655 11.375 3.195 ;
        RECT  11.115 0.655 11.165 1.255 ;
        RECT  11.115 2.255 11.165 3.195 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.580 0.880 6.775 1.200 ;
        RECT  6.580 2.165 6.625 2.765 ;
        RECT  6.565 0.880 6.580 2.765 ;
        RECT  6.420 0.940 6.565 2.765 ;
        RECT  6.345 0.940 6.420 1.200 ;
        END
        ANTENNADIFFAREA     1.0901 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.455 7.695 2.345 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 1.440 5.485 1.805 ;
        RECT  5.185 1.290 5.395 1.805 ;
        RECT  5.170 1.440 5.185 1.805 ;
        END
        ANTENNAGATEAREA     1.0751 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.540 0.530 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.815 -0.250 11.500 0.250 ;
        RECT  10.655 -0.250 10.815 1.255 ;
        RECT  7.905 -0.250 10.655 0.250 ;
        RECT  7.645 -0.250 7.905 0.405 ;
        RECT  5.285 -0.250 7.645 0.250 ;
        RECT  5.025 -0.250 5.285 0.405 ;
        RECT  0.925 -0.250 5.025 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.820 3.440 11.500 3.940 ;
        RECT  10.770 3.285 10.820 3.940 ;
        RECT  10.610 2.215 10.770 3.940 ;
        RECT  10.560 3.285 10.610 3.940 ;
        RECT  7.870 3.440 10.560 3.940 ;
        RECT  7.610 2.940 7.870 3.940 ;
        RECT  5.605 3.440 7.610 3.940 ;
        RECT  5.345 3.285 5.605 3.940 ;
        RECT  1.110 3.440 5.345 3.940 ;
        RECT  0.850 2.610 1.110 3.940 ;
        RECT  0.000 3.440 0.850 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.825 1.510 10.985 2.020 ;
        RECT  10.420 1.860 10.825 2.020 ;
        RECT  10.315 0.775 10.475 1.675 ;
        RECT  10.260 1.860 10.420 3.105 ;
        RECT  9.045 0.775 10.315 0.935 ;
        RECT  9.565 2.945 10.260 3.105 ;
        RECT  10.030 2.110 10.080 2.710 ;
        RECT  9.870 1.115 10.030 2.710 ;
        RECT  9.745 1.115 9.870 1.375 ;
        RECT  9.405 1.115 9.565 3.105 ;
        RECT  8.700 0.430 9.520 0.590 ;
        RECT  9.235 1.115 9.405 1.375 ;
        RECT  9.065 1.695 9.225 2.720 ;
        RECT  6.965 2.560 9.065 2.720 ;
        RECT  8.885 0.775 9.045 1.220 ;
        RECT  8.725 0.960 8.885 2.270 ;
        RECT  8.330 0.960 8.725 1.220 ;
        RECT  8.410 2.110 8.725 2.270 ;
        RECT  8.540 0.430 8.700 0.750 ;
        RECT  8.035 0.590 8.540 0.750 ;
        RECT  8.380 1.565 8.540 1.825 ;
        RECT  8.150 2.110 8.410 2.370 ;
        RECT  8.035 1.565 8.380 1.725 ;
        RECT  7.875 0.590 8.035 1.725 ;
        RECT  7.175 0.590 7.875 0.750 ;
        RECT  7.305 0.940 7.365 1.200 ;
        RECT  7.145 0.940 7.305 2.345 ;
        RECT  7.015 0.505 7.175 0.750 ;
        RECT  7.105 0.940 7.145 1.200 ;
        RECT  6.165 0.505 7.015 0.665 ;
        RECT  6.805 1.700 6.965 3.105 ;
        RECT  6.760 1.700 6.805 1.975 ;
        RECT  4.950 2.945 6.805 3.105 ;
        RECT  6.165 1.705 6.235 1.965 ;
        RECT  6.005 0.505 6.165 1.965 ;
        RECT  5.885 2.165 6.145 2.765 ;
        RECT  4.845 0.585 6.005 0.745 ;
        RECT  5.825 2.165 5.885 2.325 ;
        RECT  5.665 0.940 5.825 2.325 ;
        RECT  5.565 0.940 5.665 1.200 ;
        RECT  4.965 2.020 5.065 2.620 ;
        RECT  4.805 1.365 4.965 2.620 ;
        RECT  4.790 2.945 4.950 3.165 ;
        RECT  4.685 0.500 4.845 0.745 ;
        RECT  4.745 1.365 4.805 1.525 ;
        RECT  2.195 3.005 4.790 3.165 ;
        RECT  4.485 0.960 4.745 1.525 ;
        RECT  4.095 0.500 4.685 0.660 ;
        RECT  4.455 2.020 4.555 2.620 ;
        RECT  3.985 1.260 4.485 1.525 ;
        RECT  4.295 1.840 4.455 2.800 ;
        RECT  3.755 1.840 4.295 2.000 ;
        RECT  2.735 2.640 4.295 2.800 ;
        RECT  3.935 0.470 4.095 0.660 ;
        RECT  3.785 2.180 4.045 2.440 ;
        RECT  3.935 1.265 3.985 1.525 ;
        RECT  3.415 0.470 3.935 0.630 ;
        RECT  3.415 2.180 3.785 2.340 ;
        RECT  3.595 0.810 3.755 2.000 ;
        RECT  3.255 0.470 3.415 2.340 ;
        RECT  3.035 0.750 3.255 1.010 ;
        RECT  2.915 1.340 3.075 2.460 ;
        RECT  2.735 1.340 2.915 1.500 ;
        RECT  2.575 0.495 2.735 1.500 ;
        RECT  2.575 1.685 2.735 2.800 ;
        RECT  1.265 0.495 2.575 0.655 ;
        RECT  2.395 1.685 2.575 1.845 ;
        RECT  2.235 0.835 2.395 1.845 ;
        RECT  1.605 0.835 2.235 0.995 ;
        RECT  2.055 2.335 2.195 3.165 ;
        RECT  2.030 1.175 2.055 3.165 ;
        RECT  1.895 1.175 2.030 2.935 ;
        RECT  1.605 2.175 1.685 3.115 ;
        RECT  1.445 0.835 1.605 3.115 ;
        RECT  1.305 1.025 1.445 1.285 ;
        RECT  1.425 2.175 1.445 3.115 ;
        RECT  1.105 0.495 1.265 0.755 ;
        RECT  1.015 1.470 1.215 1.730 ;
        RECT  0.385 0.595 1.105 0.755 ;
        RECT  0.855 1.035 1.015 2.330 ;
        RECT  0.385 1.035 0.855 1.195 ;
        RECT  0.560 2.170 0.855 2.330 ;
        RECT  0.300 2.170 0.560 3.110 ;
        RECT  0.125 0.595 0.385 1.195 ;
    END
END AFHCONX2

MACRO AFHCINX4
    CLASS CORE ;
    FOREIGN AFHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.970 0.925 10.245 1.085 ;
        RECT  9.970 1.290 9.995 2.110 ;
        RECT  9.810 0.925 9.970 2.595 ;
        RECT  9.645 0.925 9.810 1.085 ;
        RECT  9.785 1.290 9.810 2.110 ;
        RECT  9.785 2.400 9.810 2.595 ;
        RECT  9.345 2.435 9.785 2.595 ;
        RECT  9.185 2.435 9.345 2.825 ;
        END
        ANTENNADIFFAREA     0.5288 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.335 0.810 8.495 1.240 ;
        RECT  7.475 0.810 8.335 0.970 ;
        RECT  7.555 2.745 7.715 3.220 ;
        RECT  6.775 3.060 7.555 3.220 ;
        RECT  7.315 0.810 7.475 1.765 ;
        RECT  6.775 1.605 7.315 1.765 ;
        RECT  6.535 1.605 6.775 3.220 ;
        END
        ANTENNADIFFAREA     1.3635 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.135 1.515 14.205 1.775 ;
        RECT  13.925 1.515 14.135 1.990 ;
        RECT  13.605 1.515 13.925 1.775 ;
        END
        ANTENNAGATEAREA     1.1024 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 1.700 5.575 2.025 ;
        END
        ANTENNAGATEAREA     0.7865 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.380 1.500 0.440 1.760 ;
        RECT  0.230 1.500 0.380 1.990 ;
        RECT  0.150 1.550 0.230 1.990 ;
        RECT  0.125 1.700 0.150 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.055 -0.250 15.180 0.250 ;
        RECT  14.795 -0.250 15.055 1.095 ;
        RECT  14.035 -0.250 14.795 0.250 ;
        RECT  13.775 -0.250 14.035 1.095 ;
        RECT  12.965 -0.250 13.775 0.250 ;
        RECT  12.805 -0.250 12.965 1.095 ;
        RECT  10.145 -0.250 12.805 0.250 ;
        RECT  9.545 -0.250 10.145 0.405 ;
        RECT  5.895 -0.250 9.545 0.250 ;
        RECT  5.635 -0.250 5.895 0.405 ;
        RECT  0.925 -0.250 5.635 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.055 3.440 15.180 3.940 ;
        RECT  14.795 2.105 15.055 3.940 ;
        RECT  13.995 3.440 14.795 3.940 ;
        RECT  13.735 2.895 13.995 3.940 ;
        RECT  12.875 3.440 13.735 3.940 ;
        RECT  12.685 3.285 12.875 3.940 ;
        RECT  12.465 2.895 12.685 3.940 ;
        RECT  12.275 3.285 12.465 3.940 ;
        RECT  9.905 3.440 12.275 3.940 ;
        RECT  9.645 2.785 9.905 3.940 ;
        RECT  8.835 3.440 9.645 3.940 ;
        RECT  8.675 2.565 8.835 3.940 ;
        RECT  5.685 3.440 8.675 3.940 ;
        RECT  5.405 2.205 5.685 3.940 ;
        RECT  0.905 3.440 5.405 3.940 ;
        RECT  0.645 2.530 0.905 3.940 ;
        RECT  0.000 3.440 0.645 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.385 0.595 14.545 3.110 ;
        RECT  14.285 0.595 14.385 1.195 ;
        RECT  14.285 2.170 14.385 3.110 ;
        RECT  12.625 2.395 14.285 2.555 ;
        RECT  13.425 0.595 13.525 1.195 ;
        RECT  13.425 1.955 13.445 2.215 ;
        RECT  13.265 0.595 13.425 2.215 ;
        RECT  13.185 1.275 13.265 2.215 ;
        RECT  12.625 1.275 13.185 1.435 ;
        RECT  12.465 0.470 12.625 1.435 ;
        RECT  12.465 1.615 12.625 2.555 ;
        RECT  10.485 0.470 12.465 0.630 ;
        RECT  12.285 2.395 12.465 2.555 ;
        RECT  12.125 1.035 12.285 1.455 ;
        RECT  12.125 2.395 12.285 2.905 ;
        RECT  11.945 1.295 12.125 1.455 ;
        RECT  10.895 2.745 12.125 2.905 ;
        RECT  11.785 1.295 11.945 2.565 ;
        RECT  11.605 0.855 11.825 1.115 ;
        RECT  11.755 2.305 11.785 2.565 ;
        RECT  11.445 0.810 11.605 2.105 ;
        RECT  10.825 0.810 11.445 0.970 ;
        RECT  11.405 1.945 11.445 2.105 ;
        RECT  11.245 1.945 11.405 2.565 ;
        RECT  11.165 1.150 11.265 1.310 ;
        RECT  11.005 1.150 11.165 1.765 ;
        RECT  10.895 1.605 11.005 1.765 ;
        RECT  10.735 1.605 10.895 2.905 ;
        RECT  10.665 0.810 10.825 1.425 ;
        RECT  10.515 0.970 10.665 1.425 ;
        RECT  10.385 1.265 10.515 1.425 ;
        RECT  10.325 0.470 10.485 0.745 ;
        RECT  10.225 1.265 10.385 3.205 ;
        RECT  9.175 0.585 10.325 0.745 ;
        RECT  10.085 2.945 10.225 3.205 ;
        RECT  9.445 1.345 9.605 2.255 ;
        RECT  9.175 1.345 9.445 1.505 ;
        RECT  8.495 2.095 9.445 2.255 ;
        RECT  8.835 1.755 9.265 1.915 ;
        RECT  9.015 0.585 9.175 1.505 ;
        RECT  8.675 0.470 8.835 1.915 ;
        RECT  7.085 0.470 8.675 0.630 ;
        RECT  8.155 1.755 8.675 1.915 ;
        RECT  8.335 2.095 8.495 2.440 ;
        RECT  8.225 2.280 8.335 2.440 ;
        RECT  8.065 2.280 8.225 2.920 ;
        RECT  7.995 1.755 8.155 2.090 ;
        RECT  7.815 2.280 8.065 2.440 ;
        RECT  7.815 1.150 8.035 1.310 ;
        RECT  7.655 1.150 7.815 2.440 ;
        RECT  7.205 2.280 7.655 2.440 ;
        RECT  7.045 2.280 7.205 2.880 ;
        RECT  6.925 0.470 7.085 1.085 ;
        RECT  6.355 1.265 7.015 1.425 ;
        RECT  4.905 0.925 6.925 1.085 ;
        RECT  6.245 0.430 6.710 0.590 ;
        RECT  6.225 1.265 6.355 2.365 ;
        RECT  6.085 0.430 6.245 0.745 ;
        RECT  6.195 1.265 6.225 3.145 ;
        RECT  6.175 1.265 6.195 1.425 ;
        RECT  5.965 2.205 6.195 3.145 ;
        RECT  5.245 0.585 6.085 0.745 ;
        RECT  5.915 1.610 6.015 1.870 ;
        RECT  5.755 1.265 5.915 1.870 ;
        RECT  4.935 1.265 5.755 1.425 ;
        RECT  5.085 0.470 5.245 0.745 ;
        RECT  4.935 2.205 5.125 3.145 ;
        RECT  3.885 0.470 5.085 0.630 ;
        RECT  4.865 1.265 4.935 3.145 ;
        RECT  4.745 0.810 4.905 1.085 ;
        RECT  4.775 1.265 4.865 2.365 ;
        RECT  4.225 0.810 4.745 0.970 ;
        RECT  4.405 1.150 4.565 3.220 ;
        RECT  1.415 3.060 4.405 3.220 ;
        RECT  4.065 0.810 4.225 2.880 ;
        RECT  2.975 2.720 4.065 2.880 ;
        RECT  3.725 0.470 3.885 2.510 ;
        RECT  3.265 0.745 3.425 2.335 ;
        RECT  3.255 0.745 3.265 1.005 ;
        RECT  3.165 1.750 3.265 2.335 ;
        RECT  3.095 0.485 3.255 1.005 ;
        RECT  2.435 1.750 3.165 1.910 ;
        RECT  2.375 0.485 3.095 0.645 ;
        RECT  2.715 2.585 2.975 2.880 ;
        RECT  2.655 0.855 2.915 1.035 ;
        RECT  1.925 2.720 2.715 2.880 ;
        RECT  1.975 0.875 2.655 1.035 ;
        RECT  2.275 1.750 2.435 2.495 ;
        RECT  2.115 0.435 2.375 0.695 ;
        RECT  2.175 2.235 2.275 2.495 ;
        RECT  1.470 0.485 2.115 0.645 ;
        RECT  1.925 0.875 1.975 1.205 ;
        RECT  1.765 0.875 1.925 2.880 ;
        RECT  1.715 0.875 1.765 1.205 ;
        RECT  1.665 2.150 1.765 2.880 ;
        RECT  1.310 0.485 1.470 0.845 ;
        RECT  1.415 1.035 1.465 1.295 ;
        RECT  1.255 1.035 1.415 3.220 ;
        RECT  0.945 0.685 1.310 0.845 ;
        RECT  1.205 1.035 1.255 1.295 ;
        RECT  1.155 2.185 1.255 3.220 ;
        RECT  0.945 1.500 1.045 1.760 ;
        RECT  0.785 0.685 0.945 2.330 ;
        RECT  0.385 1.035 0.785 1.195 ;
        RECT  0.395 2.170 0.785 2.330 ;
        RECT  0.135 2.170 0.395 3.110 ;
        RECT  0.125 0.595 0.385 1.195 ;
    END
END AFHCINX4

MACRO AFHCINX2
    CLASS CORE ;
    FOREIGN AFHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.340 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.615 0.925 9.175 1.085 ;
        RECT  8.590 2.395 8.645 2.995 ;
        RECT  8.590 0.925 8.615 2.110 ;
        RECT  8.430 0.925 8.590 2.995 ;
        RECT  8.405 1.290 8.430 2.110 ;
        RECT  8.385 2.395 8.430 2.995 ;
        END
        ANTENNADIFFAREA     0.5372 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.525 2.875 7.685 3.165 ;
        RECT  6.775 2.875 7.525 3.035 ;
        RECT  7.355 0.810 7.475 1.425 ;
        RECT  7.315 0.810 7.355 1.765 ;
        RECT  7.195 1.265 7.315 1.765 ;
        RECT  6.775 1.605 7.195 1.765 ;
        RECT  6.615 1.605 6.775 3.035 ;
        RECT  6.565 1.605 6.615 2.810 ;
        RECT  6.475 1.605 6.565 2.805 ;
        END
        ANTENNADIFFAREA     1.0220 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.005 1.290 13.215 1.775 ;
        RECT  12.835 1.515 13.005 1.775 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 1.700 5.565 2.025 ;
        END
        ANTENNAGATEAREA     0.7865 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.380 1.500 0.440 1.760 ;
        RECT  0.230 1.500 0.380 1.990 ;
        RECT  0.150 1.550 0.230 1.990 ;
        RECT  0.125 1.700 0.150 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.215 -0.250 13.340 0.250 ;
        RECT  12.955 -0.250 13.215 1.095 ;
        RECT  11.655 -0.250 12.955 0.250 ;
        RECT  11.395 -0.250 11.655 0.405 ;
        RECT  8.905 -0.250 11.395 0.250 ;
        RECT  8.645 -0.250 8.905 0.405 ;
        RECT  5.895 -0.250 8.645 0.250 ;
        RECT  5.635 -0.250 5.895 0.405 ;
        RECT  0.925 -0.250 5.635 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.215 3.440 13.340 3.940 ;
        RECT  12.955 2.105 13.215 3.940 ;
        RECT  11.655 3.440 12.955 3.940 ;
        RECT  11.395 3.285 11.655 3.940 ;
        RECT  9.185 3.440 11.395 3.940 ;
        RECT  8.925 2.970 9.185 3.940 ;
        RECT  8.135 3.440 8.925 3.940 ;
        RECT  7.875 2.445 8.135 3.940 ;
        RECT  5.660 3.440 7.875 3.940 ;
        RECT  5.380 2.205 5.660 3.940 ;
        RECT  0.905 3.440 5.380 3.940 ;
        RECT  0.645 2.530 0.905 3.940 ;
        RECT  0.000 3.440 0.645 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.655 0.595 12.705 1.195 ;
        RECT  12.655 2.170 12.705 3.110 ;
        RECT  12.495 0.595 12.655 3.110 ;
        RECT  12.445 0.595 12.495 1.195 ;
        RECT  12.445 2.170 12.495 3.110 ;
        RECT  11.495 2.735 12.445 2.895 ;
        RECT  12.145 0.595 12.195 1.195 ;
        RECT  12.145 1.955 12.195 2.555 ;
        RECT  11.985 0.585 12.145 2.555 ;
        RECT  11.935 0.585 11.985 1.195 ;
        RECT  11.935 1.955 11.985 2.555 ;
        RECT  11.145 0.585 11.935 0.745 ;
        RECT  11.335 1.475 11.495 3.105 ;
        RECT  10.045 2.945 11.335 3.105 ;
        RECT  10.985 0.470 11.145 0.745 ;
        RECT  11.065 2.430 11.115 2.690 ;
        RECT  10.905 1.035 11.065 2.690 ;
        RECT  9.265 0.470 10.985 0.630 ;
        RECT  10.855 2.430 10.905 2.690 ;
        RECT  10.555 0.950 10.605 1.210 ;
        RECT  10.505 0.950 10.555 2.720 ;
        RECT  10.395 0.810 10.505 2.720 ;
        RECT  10.345 0.810 10.395 1.210 ;
        RECT  9.605 0.810 10.345 0.970 ;
        RECT  9.885 1.150 10.045 3.105 ;
        RECT  9.785 1.150 9.885 1.310 ;
        RECT  9.535 0.810 9.605 1.465 ;
        RECT  9.445 0.810 9.535 2.720 ;
        RECT  9.375 1.305 9.445 2.720 ;
        RECT  9.235 2.090 9.375 2.350 ;
        RECT  9.105 0.470 9.265 0.745 ;
        RECT  8.155 0.585 9.105 0.745 ;
        RECT  7.995 0.585 8.155 2.255 ;
        RECT  7.145 2.095 7.995 2.255 ;
        RECT  7.655 0.470 7.815 1.915 ;
        RECT  7.085 0.470 7.655 0.630 ;
        RECT  7.555 1.755 7.655 1.915 ;
        RECT  6.985 2.095 7.145 2.695 ;
        RECT  6.925 0.470 7.085 1.085 ;
        RECT  6.295 1.265 7.015 1.425 ;
        RECT  4.905 0.925 6.925 1.085 ;
        RECT  6.235 0.430 6.710 0.590 ;
        RECT  6.175 1.265 6.295 2.365 ;
        RECT  6.075 0.430 6.235 0.745 ;
        RECT  6.135 1.265 6.175 3.145 ;
        RECT  5.915 2.205 6.135 3.145 ;
        RECT  5.245 0.585 6.075 0.745 ;
        RECT  5.795 1.265 5.955 1.870 ;
        RECT  4.935 1.265 5.795 1.425 ;
        RECT  5.085 0.470 5.245 0.745 ;
        RECT  4.935 2.205 5.125 3.145 ;
        RECT  3.885 0.470 5.085 0.630 ;
        RECT  4.865 1.265 4.935 3.145 ;
        RECT  4.745 0.810 4.905 1.085 ;
        RECT  4.775 1.265 4.865 2.365 ;
        RECT  4.225 0.810 4.745 0.970 ;
        RECT  4.405 1.150 4.565 3.220 ;
        RECT  1.415 3.060 4.405 3.220 ;
        RECT  4.065 0.810 4.225 2.880 ;
        RECT  2.975 2.720 4.065 2.880 ;
        RECT  3.725 0.470 3.885 2.510 ;
        RECT  3.265 0.745 3.425 2.335 ;
        RECT  3.255 0.745 3.265 1.005 ;
        RECT  3.165 1.750 3.265 2.335 ;
        RECT  3.095 0.485 3.255 1.005 ;
        RECT  2.435 1.750 3.165 1.910 ;
        RECT  2.375 0.485 3.095 0.645 ;
        RECT  2.715 2.585 2.975 2.880 ;
        RECT  2.655 0.855 2.915 1.035 ;
        RECT  1.925 2.720 2.715 2.880 ;
        RECT  1.975 0.875 2.655 1.035 ;
        RECT  2.275 1.750 2.435 2.495 ;
        RECT  2.115 0.435 2.375 0.695 ;
        RECT  2.175 2.235 2.275 2.495 ;
        RECT  1.470 0.485 2.115 0.645 ;
        RECT  1.925 0.875 1.975 1.205 ;
        RECT  1.765 0.875 1.925 2.880 ;
        RECT  1.715 0.875 1.765 1.205 ;
        RECT  1.665 2.150 1.765 2.880 ;
        RECT  1.310 0.485 1.470 0.845 ;
        RECT  1.415 1.035 1.465 1.295 ;
        RECT  1.255 1.035 1.415 3.220 ;
        RECT  0.945 0.685 1.310 0.845 ;
        RECT  1.205 1.035 1.255 1.295 ;
        RECT  1.155 2.185 1.255 3.220 ;
        RECT  0.945 1.500 1.045 1.760 ;
        RECT  0.785 0.685 0.945 2.330 ;
        RECT  0.385 1.035 0.785 1.195 ;
        RECT  0.395 2.170 0.785 2.330 ;
        RECT  0.135 2.170 0.395 3.110 ;
        RECT  0.125 0.595 0.385 1.195 ;
    END
END AFHCINX2

MACRO CMPR32X4
    CLASS CORE ;
    FOREIGN CMPR32X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.995 1.520 10.000 2.405 ;
        RECT  9.945 0.920 9.995 2.585 ;
        RECT  9.940 0.920 9.945 2.990 ;
        RECT  9.760 0.610 9.940 2.990 ;
        RECT  9.755 0.610 9.760 1.760 ;
        RECT  9.685 2.050 9.760 2.990 ;
        RECT  9.680 0.610 9.755 1.210 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.905 1.925 8.925 2.300 ;
        RECT  8.900 0.545 8.920 1.145 ;
        RECT  8.900 1.520 8.905 2.300 ;
        RECT  8.665 0.545 8.900 2.300 ;
        RECT  8.660 0.545 8.665 1.990 ;
        RECT  8.405 1.290 8.660 1.990 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 1.310 6.365 1.570 ;
        RECT  6.315 2.260 6.320 2.520 ;
        RECT  6.105 1.310 6.315 2.520 ;
        RECT  6.060 2.260 6.105 2.520 ;
        END
        ANTENNAGATEAREA     0.1976 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.490 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.510 3.165 1.990 ;
        RECT  2.645 1.510 2.885 1.825 ;
        END
        ANTENNAGATEAREA     0.2730 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.450 -0.250 10.580 0.250 ;
        RECT  10.190 -0.250 10.450 1.210 ;
        RECT  9.430 -0.250 10.190 0.250 ;
        RECT  9.170 -0.250 9.430 1.185 ;
        RECT  8.410 -0.250 9.170 0.250 ;
        RECT  8.150 -0.250 8.410 1.095 ;
        RECT  6.480 -0.250 8.150 0.250 ;
        RECT  6.220 -0.250 6.480 0.405 ;
        RECT  3.115 -0.250 6.220 0.250 ;
        RECT  2.855 -0.250 3.115 0.585 ;
        RECT  0.925 -0.250 2.855 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.455 3.440 10.580 3.940 ;
        RECT  10.195 2.140 10.455 3.940 ;
        RECT  9.435 3.440 10.195 3.940 ;
        RECT  9.175 2.920 9.435 3.940 ;
        RECT  8.385 3.440 9.175 3.940 ;
        RECT  8.125 3.285 8.385 3.940 ;
        RECT  6.420 3.440 8.125 3.940 ;
        RECT  6.160 3.285 6.420 3.940 ;
        RECT  3.155 3.440 6.160 3.940 ;
        RECT  2.895 3.285 3.155 3.940 ;
        RECT  0.925 3.440 2.895 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.475 1.510 9.575 1.770 ;
        RECT  9.315 1.510 9.475 2.735 ;
        RECT  7.330 2.575 9.315 2.735 ;
        RECT  6.760 2.915 8.075 3.075 ;
        RECT  7.800 1.035 7.900 1.295 ;
        RECT  7.800 2.135 7.870 2.395 ;
        RECT  7.640 0.595 7.800 2.395 ;
        RECT  5.935 0.595 7.640 0.755 ;
        RECT  7.610 2.135 7.640 2.395 ;
        RECT  7.290 1.035 7.390 1.295 ;
        RECT  7.290 2.280 7.330 2.735 ;
        RECT  7.170 1.035 7.290 2.735 ;
        RECT  7.130 1.035 7.170 2.540 ;
        RECT  7.070 2.280 7.130 2.540 ;
        RECT  6.720 1.035 6.880 1.295 ;
        RECT  6.720 2.145 6.820 2.405 ;
        RECT  6.600 2.735 6.760 3.075 ;
        RECT  6.560 0.935 6.720 2.405 ;
        RECT  5.450 2.735 6.600 2.895 ;
        RECT  5.550 0.935 6.560 1.095 ;
        RECT  5.775 0.485 5.935 0.755 ;
        RECT  5.790 1.275 5.890 1.435 ;
        RECT  5.630 1.275 5.790 2.545 ;
        RECT  4.050 0.485 5.775 0.645 ;
        RECT  5.250 0.825 5.550 1.095 ;
        RECT  5.290 1.275 5.450 2.895 ;
        RECT  5.120 1.275 5.290 1.435 ;
        RECT  4.810 2.735 5.290 2.895 ;
        RECT  4.480 0.825 5.250 0.985 ;
        RECT  4.950 1.615 5.110 2.555 ;
        RECT  4.820 1.615 4.950 1.775 ;
        RECT  4.560 2.395 4.950 2.555 ;
        RECT  4.660 1.225 4.820 1.775 ;
        RECT  4.480 1.955 4.770 2.215 ;
        RECT  4.460 2.395 4.560 2.795 ;
        RECT  4.320 0.825 4.480 2.215 ;
        RECT  4.400 2.395 4.460 3.015 ;
        RECT  4.300 2.535 4.400 3.015 ;
        RECT  4.050 2.055 4.320 2.215 ;
        RECT  3.710 2.855 4.300 3.015 ;
        RECT  3.540 1.520 4.140 1.780 ;
        RECT  3.890 0.485 4.050 1.315 ;
        RECT  3.950 2.055 4.050 2.425 ;
        RECT  3.840 2.055 3.950 2.670 ;
        RECT  3.790 0.765 3.890 1.315 ;
        RECT  3.790 2.165 3.840 2.670 ;
        RECT  2.530 0.765 3.790 0.925 ;
        RECT  2.320 2.510 3.790 2.670 ;
        RECT  3.450 2.855 3.710 3.115 ;
        RECT  3.380 1.105 3.540 2.330 ;
        RECT  2.320 2.855 3.450 3.015 ;
        RECT  2.305 1.105 3.380 1.265 ;
        RECT  2.660 2.170 3.380 2.330 ;
        RECT  2.500 2.035 2.660 2.330 ;
        RECT  2.370 0.685 2.530 0.925 ;
        RECT  2.355 2.035 2.500 2.195 ;
        RECT  1.665 0.685 2.370 0.845 ;
        RECT  2.175 2.395 2.320 2.670 ;
        RECT  2.160 2.855 2.320 3.260 ;
        RECT  2.160 1.595 2.175 2.670 ;
        RECT  2.015 1.595 2.160 2.555 ;
        RECT  1.495 3.100 2.160 3.260 ;
        RECT  2.005 1.595 2.015 1.755 ;
        RECT  1.845 1.055 2.005 1.755 ;
        RECT  1.835 2.760 1.980 2.920 ;
        RECT  1.665 2.025 1.835 2.285 ;
        RECT  1.675 2.540 1.835 2.920 ;
        RECT  1.325 2.540 1.675 2.700 ;
        RECT  1.505 0.685 1.665 2.285 ;
        RECT  1.335 2.945 1.495 3.260 ;
        RECT  0.385 2.945 1.335 3.105 ;
        RECT  1.165 0.975 1.325 2.700 ;
        RECT  1.075 0.975 1.165 1.235 ;
        RECT  1.065 1.990 1.165 2.700 ;
        RECT  0.745 1.500 0.985 1.760 ;
        RECT  0.585 1.135 0.745 2.330 ;
        RECT  0.385 1.135 0.585 1.295 ;
        RECT  0.385 2.170 0.585 2.330 ;
        RECT  0.125 0.600 0.385 1.295 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END CMPR32X4

MACRO CMPR32X2
    CLASS CORE ;
    FOREIGN CMPR32X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.325 0.695 9.535 2.945 ;
        RECT  9.275 0.695 9.325 1.295 ;
        RECT  9.275 2.005 9.325 2.945 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.455 1.515 8.615 1.990 ;
        RECT  8.450 1.135 8.455 2.265 ;
        RECT  8.295 0.695 8.450 2.265 ;
        RECT  8.190 0.695 8.295 1.295 ;
        RECT  8.195 2.005 8.295 2.265 ;
        END
        ANTENNADIFFAREA     0.7195 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 2.260 6.320 2.520 ;
        RECT  6.265 1.515 6.315 2.520 ;
        RECT  6.105 1.310 6.265 2.520 ;
        RECT  6.100 1.310 6.105 1.925 ;
        RECT  6.060 2.260 6.105 2.520 ;
        END
        ANTENNAGATEAREA     0.1976 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.490 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.510 3.165 1.990 ;
        RECT  2.645 1.510 2.885 1.825 ;
        END
        ANTENNAGATEAREA     0.2704 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.995 -0.250 9.660 0.250 ;
        RECT  8.735 -0.250 8.995 1.145 ;
        RECT  6.485 -0.250 8.735 0.250 ;
        RECT  6.225 -0.250 6.485 0.405 ;
        RECT  3.115 -0.250 6.225 0.250 ;
        RECT  2.855 -0.250 3.115 0.585 ;
        RECT  0.925 -0.250 2.855 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.995 3.440 9.660 3.940 ;
        RECT  8.735 2.880 8.995 3.940 ;
        RECT  6.420 3.440 8.735 3.940 ;
        RECT  6.160 3.285 6.420 3.940 ;
        RECT  3.155 3.440 6.160 3.940 ;
        RECT  2.895 3.285 3.155 3.940 ;
        RECT  0.925 3.440 2.895 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.045 1.565 9.145 1.825 ;
        RECT  8.885 1.565 9.045 2.690 ;
        RECT  7.330 2.530 8.885 2.690 ;
        RECT  7.825 2.870 8.085 3.130 ;
        RECT  7.820 1.035 7.940 1.295 ;
        RECT  7.820 2.090 7.870 2.350 ;
        RECT  6.760 2.870 7.825 3.030 ;
        RECT  7.660 0.595 7.820 2.350 ;
        RECT  5.935 0.595 7.660 0.755 ;
        RECT  7.610 2.090 7.660 2.350 ;
        RECT  7.330 1.035 7.430 1.295 ;
        RECT  7.170 1.035 7.330 2.690 ;
        RECT  7.160 2.280 7.170 2.690 ;
        RECT  7.070 2.280 7.160 2.540 ;
        RECT  6.720 1.035 6.920 1.295 ;
        RECT  6.720 2.145 6.820 2.405 ;
        RECT  6.600 2.735 6.760 3.030 ;
        RECT  6.560 0.935 6.720 2.405 ;
        RECT  5.450 2.735 6.600 2.895 ;
        RECT  5.550 0.935 6.560 1.095 ;
        RECT  5.775 0.485 5.935 0.755 ;
        RECT  5.790 1.275 5.895 1.435 ;
        RECT  5.630 1.275 5.790 2.545 ;
        RECT  4.050 0.485 5.775 0.645 ;
        RECT  5.290 0.830 5.550 1.095 ;
        RECT  5.290 1.275 5.450 2.895 ;
        RECT  4.480 0.880 5.290 1.040 ;
        RECT  5.120 1.275 5.290 1.435 ;
        RECT  4.810 2.735 5.290 2.895 ;
        RECT  4.950 1.615 5.110 2.555 ;
        RECT  4.820 1.615 4.950 1.775 ;
        RECT  4.560 2.395 4.950 2.555 ;
        RECT  4.660 1.225 4.820 1.775 ;
        RECT  4.480 1.955 4.770 2.215 ;
        RECT  4.460 2.395 4.560 2.795 ;
        RECT  4.320 0.880 4.480 2.215 ;
        RECT  4.400 2.395 4.460 3.010 ;
        RECT  4.300 2.535 4.400 3.010 ;
        RECT  4.050 2.055 4.320 2.215 ;
        RECT  2.320 2.850 4.300 3.010 ;
        RECT  3.540 1.520 4.140 1.780 ;
        RECT  3.890 0.485 4.050 1.315 ;
        RECT  3.950 2.055 4.050 2.425 ;
        RECT  3.840 2.055 3.950 2.670 ;
        RECT  3.790 0.765 3.890 1.315 ;
        RECT  3.790 2.165 3.840 2.670 ;
        RECT  2.530 0.765 3.790 0.925 ;
        RECT  2.320 2.510 3.790 2.670 ;
        RECT  3.380 1.105 3.540 2.330 ;
        RECT  2.305 1.105 3.380 1.265 ;
        RECT  2.660 2.170 3.380 2.330 ;
        RECT  2.500 2.035 2.660 2.330 ;
        RECT  2.370 0.685 2.530 0.925 ;
        RECT  2.355 2.035 2.500 2.195 ;
        RECT  1.665 0.685 2.370 0.845 ;
        RECT  2.175 2.420 2.320 2.670 ;
        RECT  2.160 2.850 2.320 3.260 ;
        RECT  2.160 1.595 2.175 2.670 ;
        RECT  2.015 1.595 2.160 2.580 ;
        RECT  1.495 3.100 2.160 3.260 ;
        RECT  2.005 1.595 2.015 1.755 ;
        RECT  1.845 1.055 2.005 1.755 ;
        RECT  1.835 2.760 1.980 2.920 ;
        RECT  1.665 2.025 1.835 2.285 ;
        RECT  1.675 2.540 1.835 2.920 ;
        RECT  1.325 2.540 1.675 2.700 ;
        RECT  1.505 0.685 1.665 2.285 ;
        RECT  1.335 2.945 1.495 3.260 ;
        RECT  0.385 2.945 1.335 3.105 ;
        RECT  1.165 1.035 1.325 2.700 ;
        RECT  1.075 1.035 1.165 1.295 ;
        RECT  1.065 1.990 1.165 2.700 ;
        RECT  0.745 1.500 0.985 1.760 ;
        RECT  0.585 1.135 0.745 2.330 ;
        RECT  0.385 1.135 0.585 1.295 ;
        RECT  0.385 2.170 0.585 2.330 ;
        RECT  0.125 0.695 0.385 1.295 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END CMPR32X2

MACRO CMPR22X4
    CLASS CORE ;
    FOREIGN CMPR22X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.800 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.130 0.475 8.480 0.760 ;
        RECT  7.460 0.600 8.130 0.760 ;
        RECT  7.590 2.035 7.850 2.700 ;
        RECT  6.830 2.035 7.590 2.195 ;
        RECT  7.200 0.600 7.460 0.870 ;
        RECT  6.440 0.600 7.200 0.760 ;
        RECT  6.775 2.035 6.830 2.725 ;
        RECT  6.565 2.035 6.775 2.810 ;
        RECT  5.805 2.175 6.565 2.415 ;
        RECT  6.420 0.600 6.440 1.200 ;
        RECT  6.180 0.600 6.420 1.500 ;
        RECT  5.420 1.260 6.180 1.500 ;
        RECT  5.370 2.135 5.805 2.415 ;
        RECT  5.160 1.015 5.420 1.500 ;
        RECT  4.785 2.175 5.370 2.415 ;
        RECT  4.395 1.260 5.160 1.500 ;
        RECT  4.450 2.135 4.785 2.415 ;
        RECT  3.830 2.175 4.450 2.415 ;
        RECT  4.140 1.015 4.395 1.500 ;
        RECT  4.135 1.015 4.140 1.425 ;
        RECT  3.260 1.265 4.135 1.425 ;
        RECT  3.370 2.115 3.830 2.415 ;
        RECT  3.260 2.110 3.370 2.415 ;
        RECT  3.020 1.265 3.260 2.415 ;
        END
        ANTENNADIFFAREA     3.7667 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.435 0.915 13.675 2.435 ;
        RECT  13.215 0.915 13.435 1.075 ;
        RECT  13.215 2.275 13.435 2.435 ;
        RECT  13.165 0.695 13.215 1.075 ;
        RECT  13.155 2.275 13.215 2.995 ;
        RECT  12.905 0.475 13.165 1.075 ;
        RECT  12.895 2.275 13.155 3.215 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 1.430 7.995 1.690 ;
        RECT  7.735 1.430 7.945 1.840 ;
        RECT  6.315 1.680 7.735 1.840 ;
        RECT  6.130 1.680 6.315 1.990 ;
        RECT  6.105 1.700 6.130 1.990 ;
        RECT  3.705 1.715 6.105 1.875 ;
        RECT  3.445 1.625 3.705 1.875 ;
        END
        ANTENNAGATEAREA     1.7420 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.535 1.620 11.285 1.780 ;
        RECT  9.325 1.290 9.535 1.780 ;
        END
        ANTENNAGATEAREA     1.6952 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.675 -0.250 13.800 0.250 ;
        RECT  13.415 -0.250 13.675 0.735 ;
        RECT  12.655 -0.250 13.415 0.250 ;
        RECT  12.395 -0.250 12.655 0.735 ;
        RECT  11.745 -0.250 12.395 0.250 ;
        RECT  11.485 -0.250 11.745 1.075 ;
        RECT  10.725 -0.250 11.485 0.250 ;
        RECT  10.465 -0.250 10.725 1.075 ;
        RECT  9.705 -0.250 10.465 0.250 ;
        RECT  9.445 -0.250 9.705 1.075 ;
        RECT  3.655 -0.250 9.445 0.250 ;
        RECT  3.395 -0.250 3.655 0.405 ;
        RECT  2.465 -0.250 3.395 0.250 ;
        RECT  2.205 -0.250 2.465 0.405 ;
        RECT  1.405 -0.250 2.205 0.250 ;
        RECT  1.145 -0.250 1.405 1.095 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.185 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.665 3.440 13.800 3.940 ;
        RECT  13.405 2.615 13.665 3.940 ;
        RECT  12.645 3.440 13.405 3.940 ;
        RECT  12.385 2.535 12.645 3.940 ;
        RECT  11.625 3.440 12.385 3.940 ;
        RECT  11.365 2.760 11.625 3.940 ;
        RECT  10.570 3.440 11.365 3.940 ;
        RECT  10.310 2.825 10.570 3.940 ;
        RECT  9.470 3.440 10.310 3.940 ;
        RECT  9.210 3.285 9.470 3.940 ;
        RECT  8.415 3.440 9.210 3.940 ;
        RECT  8.155 3.285 8.415 3.940 ;
        RECT  3.255 3.440 8.155 3.940 ;
        RECT  2.995 3.285 3.255 3.940 ;
        RECT  2.455 3.440 2.995 3.940 ;
        RECT  2.195 3.285 2.455 3.940 ;
        RECT  1.405 3.440 2.195 3.940 ;
        RECT  1.145 2.510 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.100 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.990 1.255 13.150 2.095 ;
        RECT  12.255 1.255 12.990 1.415 ;
        RECT  12.135 1.935 12.990 2.095 ;
        RECT  11.680 1.595 12.810 1.755 ;
        RECT  11.995 1.015 12.255 1.415 ;
        RECT  11.975 1.935 12.135 3.125 ;
        RECT  11.235 1.255 11.995 1.415 ;
        RECT  11.875 2.185 11.975 3.125 ;
        RECT  11.115 2.405 11.875 2.565 ;
        RECT  11.520 1.595 11.680 2.125 ;
        RECT  8.920 1.965 11.520 2.125 ;
        RECT  10.975 0.610 11.235 1.415 ;
        RECT  10.855 2.310 11.115 2.910 ;
        RECT  10.215 1.255 10.975 1.415 ;
        RECT  10.020 2.405 10.855 2.565 ;
        RECT  10.055 0.610 10.215 1.415 ;
        RECT  9.955 0.610 10.055 1.210 ;
        RECT  9.760 2.310 10.020 2.920 ;
        RECT  8.370 2.760 9.760 2.920 ;
        RECT  8.870 1.965 8.920 2.575 ;
        RECT  8.870 1.035 8.880 1.295 ;
        RECT  8.710 1.035 8.870 2.575 ;
        RECT  8.620 1.035 8.710 1.295 ;
        RECT  8.660 1.975 8.710 2.575 ;
        RECT  8.210 1.055 8.370 3.085 ;
        RECT  7.970 1.055 8.210 1.220 ;
        RECT  7.340 2.925 8.210 3.085 ;
        RECT  7.710 0.960 7.970 1.220 ;
        RECT  6.950 1.060 7.710 1.220 ;
        RECT  7.300 2.445 7.340 3.085 ;
        RECT  7.080 2.445 7.300 3.195 ;
        RECT  6.315 3.035 7.080 3.195 ;
        RECT  6.690 0.960 6.950 1.220 ;
        RECT  6.055 2.595 6.315 3.195 ;
        RECT  2.385 2.595 6.055 2.755 ;
        RECT  5.670 0.475 5.930 1.075 ;
        RECT  4.910 0.585 5.670 0.745 ;
        RECT  5.035 2.935 5.295 3.195 ;
        RECT  4.275 2.935 5.035 3.095 ;
        RECT  4.650 0.475 4.910 1.075 ;
        RECT  1.915 0.585 4.650 0.745 ;
        RECT  4.015 2.935 4.275 3.195 ;
        RECT  1.915 2.935 4.015 3.095 ;
        RECT  2.805 0.925 3.950 1.085 ;
        RECT  2.645 0.925 2.805 2.355 ;
        RECT  2.225 1.635 2.385 2.755 ;
        RECT  1.105 1.635 2.225 1.795 ;
        RECT  1.655 0.585 1.915 1.445 ;
        RECT  1.655 2.155 1.915 3.095 ;
        RECT  0.895 1.285 1.655 1.445 ;
        RECT  0.895 2.155 1.655 2.315 ;
        RECT  0.850 0.695 0.895 1.445 ;
        RECT  0.850 2.155 0.895 3.095 ;
        RECT  0.690 0.695 0.850 3.095 ;
        RECT  0.635 0.695 0.690 1.295 ;
        RECT  0.635 2.155 0.690 3.095 ;
    END
END CMPR22X4

MACRO CMPR22X2
    CLASS CORE ;
    FOREIGN CMPR22X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.315 0.840 4.575 1.215 ;
        RECT  4.135 2.110 4.395 2.710 ;
        RECT  3.555 1.055 4.315 1.215 ;
        RECT  3.990 2.110 4.135 2.400 ;
        RECT  3.555 2.110 3.990 2.270 ;
        RECT  3.345 0.480 3.555 1.215 ;
        RECT  3.375 2.110 3.555 2.400 ;
        RECT  3.115 2.110 3.375 2.715 ;
        RECT  3.295 0.480 3.345 1.080 ;
        RECT  2.545 0.920 3.295 1.080 ;
        RECT  2.545 2.110 3.115 2.270 ;
        RECT  2.385 0.820 2.545 2.280 ;
        RECT  2.275 0.820 2.385 1.080 ;
        RECT  2.355 2.110 2.385 2.280 ;
        RECT  2.095 2.110 2.355 2.395 ;
        END
        ANTENNADIFFAREA     2.1834 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.595 0.625 8.615 3.000 ;
        RECT  8.405 0.625 8.595 3.115 ;
        RECT  8.355 0.625 8.405 1.225 ;
        RECT  8.335 2.175 8.405 3.115 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.255 1.470 4.535 1.730 ;
        RECT  3.095 1.520 4.255 1.730 ;
        RECT  2.890 1.290 3.095 1.730 ;
        RECT  2.885 1.290 2.890 1.900 ;
        RECT  2.730 1.570 2.885 1.900 ;
        END
        ANTENNAGATEAREA     0.8749 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 1.685 6.515 1.845 ;
        RECT  5.185 1.685 5.395 1.990 ;
        END
        ANTENNAGATEAREA     0.8853 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.105 -0.250 8.740 0.250 ;
        RECT  7.845 -0.250 8.105 1.075 ;
        RECT  7.045 -0.250 7.845 0.250 ;
        RECT  6.785 -0.250 7.045 0.795 ;
        RECT  5.945 -0.250 6.785 0.250 ;
        RECT  5.685 -0.250 5.945 0.765 ;
        RECT  1.445 -0.250 5.685 0.250 ;
        RECT  1.185 -0.250 1.445 0.405 ;
        RECT  0.385 -0.250 1.185 0.250 ;
        RECT  0.125 -0.250 0.385 1.195 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.085 3.440 8.740 3.940 ;
        RECT  7.825 2.460 8.085 3.940 ;
        RECT  7.065 3.440 7.825 3.940 ;
        RECT  6.805 2.835 7.065 3.940 ;
        RECT  6.005 3.440 6.805 3.940 ;
        RECT  5.745 2.945 6.005 3.940 ;
        RECT  4.905 3.440 5.745 3.940 ;
        RECT  4.645 3.285 4.905 3.940 ;
        RECT  1.445 3.440 4.645 3.940 ;
        RECT  1.185 3.285 1.445 3.940 ;
        RECT  0.385 3.440 1.185 3.940 ;
        RECT  0.125 2.935 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.955 1.255 8.115 2.265 ;
        RECT  7.595 1.255 7.955 1.415 ;
        RECT  7.575 2.105 7.955 2.265 ;
        RECT  7.610 1.600 7.770 1.860 ;
        RECT  7.055 1.650 7.610 1.810 ;
        RECT  7.435 0.600 7.595 1.415 ;
        RECT  7.315 2.105 7.575 3.045 ;
        RECT  7.335 0.600 7.435 1.200 ;
        RECT  6.495 0.995 7.335 1.155 ;
        RECT  6.555 2.450 7.315 2.610 ;
        RECT  6.895 1.345 7.055 2.250 ;
        RECT  5.085 1.345 6.895 1.505 ;
        RECT  6.020 2.090 6.895 2.250 ;
        RECT  6.295 2.450 6.555 3.150 ;
        RECT  6.235 0.555 6.495 1.155 ;
        RECT  4.785 2.595 6.295 2.755 ;
        RECT  5.470 0.995 6.235 1.155 ;
        RECT  5.860 2.090 6.020 2.405 ;
        RECT  4.985 2.245 5.860 2.405 ;
        RECT  5.310 0.500 5.470 1.155 ;
        RECT  4.065 0.500 5.310 0.660 ;
        RECT  4.985 1.005 5.085 1.505 ;
        RECT  4.825 1.005 4.985 2.405 ;
        RECT  4.625 2.595 4.785 3.090 ;
        RECT  3.885 2.930 4.625 3.090 ;
        RECT  3.805 0.500 4.065 0.850 ;
        RECT  3.625 2.605 3.885 3.205 ;
        RECT  0.915 2.935 3.625 3.095 ;
        RECT  2.785 0.480 3.045 0.740 ;
        RECT  2.605 2.485 2.865 2.745 ;
        RECT  1.800 0.480 2.785 0.640 ;
        RECT  1.405 2.585 2.605 2.745 ;
        RECT  1.995 1.260 2.205 1.520 ;
        RECT  1.845 0.935 1.995 1.520 ;
        RECT  1.735 0.935 1.845 2.215 ;
        RECT  1.640 0.480 1.800 0.750 ;
        RECT  1.685 1.360 1.735 2.215 ;
        RECT  1.585 1.955 1.685 2.215 ;
        RECT  0.895 0.590 1.640 0.750 ;
        RECT  1.245 1.130 1.405 2.745 ;
        RECT  0.895 1.130 1.245 1.290 ;
        RECT  0.635 2.115 1.245 2.375 ;
        RECT  0.450 1.585 1.065 1.845 ;
        RECT  0.755 2.590 0.915 3.095 ;
        RECT  0.635 0.590 0.895 1.290 ;
        RECT  0.450 2.590 0.755 2.750 ;
        RECT  0.290 1.585 0.450 2.750 ;
    END
END CMPR22X2

MACRO BMXIX4
    CLASS CORE ;
    FOREIGN BMXIX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.545 2.520 12.950 3.025 ;
        END
        ANTENNAGATEAREA     0.4524 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.615 1.475 9.330 1.735 ;
        RECT  8.405 1.475 8.615 1.990 ;
        RECT  8.390 1.475 8.405 1.735 ;
        END
        ANTENNAGATEAREA     0.6474 ;
    END S
    PIN PPN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.060 1.515 14.135 2.585 ;
        RECT  13.800 0.655 14.060 3.045 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END PPN
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 1.485 8.155 1.990 ;
        RECT  7.885 1.485 7.945 1.845 ;
        END
        ANTENNAGATEAREA     0.4524 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 1.255 3.055 2.485 ;
        RECT  2.635 2.325 2.895 2.485 ;
        RECT  2.625 2.325 2.635 2.585 ;
        RECT  2.465 2.325 2.625 2.770 ;
        RECT  2.425 2.610 2.465 2.770 ;
        RECT  2.165 2.610 2.425 3.220 ;
        RECT  0.795 2.610 2.165 2.770 ;
        RECT  0.725 2.520 0.795 2.810 ;
        RECT  0.625 1.715 0.725 2.810 ;
        RECT  0.585 1.615 0.625 2.810 ;
        RECT  0.565 1.615 0.585 2.770 ;
        RECT  0.465 1.615 0.565 1.875 ;
        END
        ANTENNAGATEAREA     0.4524 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.635 1.355 1.990 ;
        END
        ANTENNAGATEAREA     0.6448 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.570 -0.250 14.720 0.250 ;
        RECT  14.310 -0.250 14.570 1.195 ;
        RECT  13.520 -0.250 14.310 0.250 ;
        RECT  13.260 -0.250 13.520 0.405 ;
        RECT  9.370 -0.250 13.260 0.250 ;
        RECT  9.110 -0.250 9.370 0.405 ;
        RECT  8.270 -0.250 9.110 0.250 ;
        RECT  8.010 -0.250 8.270 0.405 ;
        RECT  1.845 -0.250 8.010 0.250 ;
        RECT  1.585 -0.250 1.845 0.755 ;
        RECT  0.785 -0.250 1.585 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.575 3.440 14.720 3.940 ;
        RECT  14.315 2.255 14.575 3.940 ;
        RECT  13.510 3.440 14.315 3.940 ;
        RECT  13.250 2.255 13.510 3.940 ;
        RECT  9.370 3.440 13.250 3.940 ;
        RECT  9.110 3.285 9.370 3.940 ;
        RECT  8.305 3.440 9.110 3.940 ;
        RECT  8.045 3.285 8.305 3.940 ;
        RECT  1.735 3.440 8.045 3.940 ;
        RECT  1.475 3.285 1.735 3.940 ;
        RECT  0.785 3.440 1.475 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.520 1.475 13.620 1.735 ;
        RECT  13.360 0.615 13.520 1.735 ;
        RECT  12.460 0.615 13.360 0.775 ;
        RECT  12.870 1.035 12.970 1.295 ;
        RECT  12.870 1.955 12.970 2.215 ;
        RECT  12.710 1.035 12.870 2.215 ;
        RECT  12.470 1.470 12.710 1.730 ;
        RECT  12.290 0.615 12.460 1.115 ;
        RECT  12.290 2.050 12.320 2.650 ;
        RECT  12.130 0.615 12.290 2.650 ;
        RECT  11.440 0.615 12.130 0.775 ;
        RECT  12.060 2.050 12.130 2.650 ;
        RECT  11.810 0.955 11.950 1.215 ;
        RECT  11.710 0.955 11.810 2.710 ;
        RECT  11.650 0.955 11.710 3.105 ;
        RECT  11.550 2.110 11.650 3.105 ;
        RECT  7.695 2.945 11.550 3.105 ;
        RECT  11.325 0.615 11.440 1.115 ;
        RECT  11.280 0.615 11.325 2.765 ;
        RECT  11.165 0.855 11.280 2.765 ;
        RECT  11.040 2.165 11.165 2.765 ;
        RECT  10.280 2.605 11.040 2.765 ;
        RECT  10.815 0.855 10.930 1.115 ;
        RECT  10.655 0.585 10.815 2.425 ;
        RECT  6.850 0.585 10.655 0.745 ;
        RECT  10.530 2.165 10.655 2.425 ;
        RECT  10.280 0.955 10.420 1.215 ;
        RECT  10.120 0.955 10.280 2.765 ;
        RECT  10.020 2.165 10.120 2.765 ;
        RECT  9.670 0.925 9.910 1.185 ;
        RECT  9.670 2.165 9.770 2.765 ;
        RECT  9.650 0.925 9.670 2.765 ;
        RECT  9.510 0.975 9.650 2.765 ;
        RECT  8.820 0.975 9.510 1.135 ;
        RECT  8.820 2.605 9.510 2.765 ;
        RECT  8.560 0.925 8.820 1.185 ;
        RECT  8.560 2.170 8.820 2.765 ;
        RECT  7.355 2.605 8.560 2.765 ;
        RECT  7.700 1.035 7.870 1.295 ;
        RECT  7.700 2.105 7.755 2.365 ;
        RECT  7.540 1.035 7.700 2.365 ;
        RECT  7.535 2.945 7.695 3.220 ;
        RECT  7.405 1.500 7.540 1.760 ;
        RECT  7.495 2.105 7.540 2.365 ;
        RECT  3.395 3.060 7.535 3.220 ;
        RECT  7.190 1.020 7.360 1.280 ;
        RECT  7.255 2.605 7.355 2.880 ;
        RECT  7.190 1.940 7.255 2.880 ;
        RECT  7.095 1.020 7.190 2.880 ;
        RECT  7.030 1.020 7.095 2.100 ;
        RECT  5.255 2.720 7.095 2.880 ;
        RECT  6.745 0.585 6.850 1.280 ;
        RECT  6.745 2.280 6.845 2.540 ;
        RECT  6.690 0.585 6.745 2.540 ;
        RECT  6.585 1.020 6.690 2.540 ;
        RECT  5.765 2.380 6.585 2.540 ;
        RECT  6.205 0.920 6.340 1.180 ;
        RECT  6.205 2.040 6.305 2.200 ;
        RECT  6.045 0.650 6.205 2.200 ;
        RECT  4.890 0.650 6.045 0.810 ;
        RECT  5.730 0.995 5.830 1.255 ;
        RECT  5.730 2.280 5.765 2.540 ;
        RECT  5.570 0.995 5.730 2.540 ;
        RECT  5.505 2.280 5.570 2.540 ;
        RECT  5.205 1.195 5.290 1.455 ;
        RECT  5.205 2.620 5.255 2.880 ;
        RECT  5.045 1.195 5.205 2.880 ;
        RECT  5.030 1.195 5.045 1.455 ;
        RECT  4.995 2.620 5.045 2.880 ;
        RECT  3.835 2.720 4.995 2.880 ;
        RECT  4.790 0.650 4.890 0.945 ;
        RECT  4.790 2.115 4.855 2.375 ;
        RECT  4.630 0.470 4.790 2.375 ;
        RECT  2.715 0.470 4.630 0.630 ;
        RECT  4.595 2.115 4.630 2.375 ;
        RECT  4.280 0.810 4.380 1.070 ;
        RECT  4.280 2.255 4.345 2.515 ;
        RECT  4.120 0.810 4.280 2.515 ;
        RECT  3.395 0.810 4.120 0.970 ;
        RECT  4.085 2.255 4.120 2.515 ;
        RECT  3.735 1.150 3.835 1.310 ;
        RECT  3.735 2.620 3.835 2.880 ;
        RECT  3.575 1.150 3.735 2.880 ;
        RECT  3.235 0.810 3.395 3.220 ;
        RECT  3.015 0.810 3.235 1.070 ;
        RECT  2.845 2.715 3.235 2.975 ;
        RECT  2.555 0.470 2.715 2.145 ;
        RECT  2.455 0.470 2.555 1.095 ;
        RECT  2.285 1.985 2.555 2.145 ;
        RECT  1.335 0.935 2.455 1.095 ;
        RECT  2.215 1.275 2.375 1.805 ;
        RECT  2.025 1.985 2.285 2.330 ;
        RECT  0.385 1.275 2.215 1.435 ;
        RECT  1.335 2.170 2.025 2.330 ;
        RECT  1.075 0.495 1.335 1.095 ;
        RECT  1.075 2.170 1.335 2.430 ;
        RECT  0.285 0.855 0.385 1.435 ;
        RECT  0.285 2.055 0.385 2.315 ;
        RECT  0.125 0.855 0.285 2.315 ;
    END
END BMXIX4

MACRO BMXIX2
    CLASS CORE ;
    FOREIGN BMXIX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.510 2.555 8.770 3.220 ;
        RECT  8.405 2.930 8.510 3.220 ;
        END
        ANTENNAGATEAREA     0.2275 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 1.290 6.775 1.785 ;
        RECT  6.475 1.440 6.565 1.785 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END S
    PIN PPN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.890 0.695 9.995 2.585 ;
        RECT  9.835 0.695 9.890 2.915 ;
        RECT  9.735 0.695 9.835 1.295 ;
        RECT  9.630 1.975 9.835 2.915 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END PPN
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.645 1.290 5.855 1.815 ;
        RECT  5.435 1.555 5.645 1.815 ;
        END
        ANTENNAGATEAREA     0.2275 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.455 1.490 2.615 2.780 ;
        RECT  2.105 2.620 2.455 2.780 ;
        RECT  2.005 2.620 2.105 2.880 ;
        RECT  1.845 2.620 2.005 3.105 ;
        RECT  0.795 2.945 1.845 3.105 ;
        RECT  0.585 1.615 0.795 3.105 ;
        RECT  0.475 1.615 0.585 1.875 ;
        END
        ANTENNAGATEAREA     0.2275 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.975 1.615 1.410 1.990 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.455 -0.250 10.120 0.250 ;
        RECT  9.195 -0.250 9.455 0.405 ;
        RECT  6.795 -0.250 9.195 0.250 ;
        RECT  5.735 -0.250 6.795 0.405 ;
        RECT  1.765 -0.250 5.735 0.250 ;
        RECT  1.505 -0.250 1.765 0.405 ;
        RECT  0.815 -0.250 1.505 0.250 ;
        RECT  0.555 -0.250 0.815 0.800 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 3.440 10.120 3.940 ;
        RECT  9.120 2.275 9.380 3.940 ;
        RECT  6.795 3.440 9.120 3.940 ;
        RECT  5.735 3.285 6.795 3.940 ;
        RECT  5.355 3.440 5.735 3.940 ;
        RECT  3.395 3.390 5.355 3.940 ;
        RECT  1.735 3.440 3.395 3.940 ;
        RECT  1.475 3.285 1.735 3.940 ;
        RECT  0.785 3.440 1.475 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.475 1.475 9.640 1.735 ;
        RECT  9.315 0.615 9.475 1.735 ;
        RECT  7.820 0.615 9.315 0.775 ;
        RECT  8.840 1.035 8.950 1.295 ;
        RECT  8.680 1.035 8.840 2.355 ;
        RECT  8.580 1.775 8.680 2.355 ;
        RECT  8.345 1.775 8.580 1.935 ;
        RECT  8.180 1.035 8.440 1.295 ;
        RECT  8.165 2.115 8.330 2.715 ;
        RECT  8.165 1.135 8.180 1.295 ;
        RECT  8.005 1.135 8.165 2.995 ;
        RECT  5.385 2.835 8.005 2.995 ;
        RECT  7.660 0.615 7.820 2.595 ;
        RECT  7.560 0.935 7.660 1.195 ;
        RECT  7.560 1.995 7.660 2.595 ;
        RECT  7.260 1.035 7.310 1.295 ;
        RECT  7.260 1.995 7.310 2.595 ;
        RECT  7.210 1.035 7.260 2.595 ;
        RECT  7.100 0.655 7.210 2.595 ;
        RECT  7.050 0.655 7.100 1.295 ;
        RECT  7.050 1.995 7.100 2.595 ;
        RECT  4.485 0.655 7.050 0.815 ;
        RECT  6.295 2.055 6.395 2.655 ;
        RECT  6.295 1.000 6.345 1.260 ;
        RECT  6.135 1.000 6.295 2.655 ;
        RECT  5.045 2.495 6.135 2.655 ;
        RECT  5.185 1.995 5.445 2.255 ;
        RECT  5.165 1.035 5.385 1.295 ;
        RECT  5.225 2.835 5.385 3.105 ;
        RECT  2.955 2.945 5.225 3.105 ;
        RECT  5.165 1.995 5.185 2.155 ;
        RECT  5.005 1.035 5.165 2.155 ;
        RECT  4.825 2.495 5.045 2.765 ;
        RECT  4.665 1.035 4.825 2.765 ;
        RECT  3.625 2.605 4.665 2.765 ;
        RECT  4.325 0.655 4.485 2.425 ;
        RECT  4.075 1.035 4.325 1.295 ;
        RECT  3.775 1.955 4.025 2.215 ;
        RECT  3.775 1.035 3.825 1.295 ;
        RECT  3.765 1.035 3.775 2.215 ;
        RECT  3.725 1.035 3.765 2.165 ;
        RECT  3.615 0.470 3.725 2.165 ;
        RECT  3.365 2.505 3.625 2.765 ;
        RECT  3.565 0.470 3.615 1.295 ;
        RECT  2.290 0.470 3.565 0.630 ;
        RECT  3.320 2.505 3.365 2.665 ;
        RECT  3.160 0.810 3.320 2.665 ;
        RECT  3.055 0.810 3.160 0.970 ;
        RECT  2.805 1.150 2.955 3.105 ;
        RECT  2.795 0.960 2.805 3.105 ;
        RECT  2.545 0.960 2.795 1.310 ;
        RECT  2.275 0.470 2.290 1.070 ;
        RECT  2.245 0.470 2.275 2.330 ;
        RECT  2.130 0.470 2.245 2.440 ;
        RECT  2.115 0.810 2.130 2.440 ;
        RECT  2.030 0.810 2.115 1.095 ;
        RECT  1.985 2.170 2.115 2.440 ;
        RECT  1.365 0.935 2.030 1.095 ;
        RECT  1.335 2.170 1.985 2.330 ;
        RECT  1.775 1.275 1.935 1.985 ;
        RECT  0.385 1.275 1.775 1.435 ;
        RECT  1.105 0.835 1.365 1.095 ;
        RECT  1.075 2.170 1.335 2.765 ;
        RECT  0.285 1.035 0.385 1.435 ;
        RECT  0.285 2.095 0.385 2.355 ;
        RECT  0.125 1.035 0.285 2.355 ;
    END
END BMXIX2

MACRO BMXX4
    CLASS CORE ;
    FOREIGN BMXX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.020 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.845 2.785 15.390 3.220 ;
        END
        ANTENNAGATEAREA     0.5902 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.615 1.475 9.330 1.735 ;
        RECT  8.405 1.475 8.615 1.990 ;
        RECT  8.390 1.475 8.405 1.735 ;
        END
        ANTENNAGATEAREA     0.6474 ;
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.380 1.105 16.435 2.585 ;
        RECT  16.120 0.655 16.380 3.045 ;
        END
        ANTENNADIFFAREA     0.8268 ;
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 1.485 8.155 1.990 ;
        RECT  7.885 1.485 7.945 1.845 ;
        END
        ANTENNAGATEAREA     0.4524 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 1.255 3.055 2.485 ;
        RECT  2.635 2.325 2.895 2.485 ;
        RECT  2.625 2.325 2.635 2.585 ;
        RECT  2.465 2.325 2.625 2.770 ;
        RECT  2.425 2.610 2.465 2.770 ;
        RECT  2.165 2.610 2.425 3.220 ;
        RECT  0.795 2.610 2.165 2.770 ;
        RECT  0.725 2.520 0.795 2.810 ;
        RECT  0.625 1.715 0.725 2.810 ;
        RECT  0.585 1.615 0.625 2.810 ;
        RECT  0.565 1.615 0.585 2.770 ;
        RECT  0.465 1.615 0.565 1.875 ;
        END
        ANTENNAGATEAREA     0.4524 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.635 1.355 1.990 ;
        END
        ANTENNAGATEAREA     0.6448 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.890 -0.250 17.020 0.250 ;
        RECT  16.630 -0.250 16.890 1.195 ;
        RECT  15.830 -0.250 16.630 0.250 ;
        RECT  15.570 -0.250 15.830 0.405 ;
        RECT  12.200 -0.250 15.570 0.250 ;
        RECT  11.940 -0.250 12.200 0.405 ;
        RECT  11.400 -0.250 11.940 0.250 ;
        RECT  11.140 -0.250 11.400 0.405 ;
        RECT  10.310 -0.250 11.140 0.250 ;
        RECT  10.050 -0.250 10.310 0.405 ;
        RECT  9.370 -0.250 10.050 0.250 ;
        RECT  9.110 -0.250 9.370 0.405 ;
        RECT  8.270 -0.250 9.110 0.250 ;
        RECT  8.010 -0.250 8.270 0.405 ;
        RECT  1.845 -0.250 8.010 0.250 ;
        RECT  1.585 -0.250 1.845 0.755 ;
        RECT  0.785 -0.250 1.585 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.890 3.440 17.020 3.940 ;
        RECT  16.630 2.255 16.890 3.940 ;
        RECT  15.855 3.440 16.630 3.940 ;
        RECT  15.595 2.255 15.855 3.940 ;
        RECT  12.070 3.440 15.595 3.940 ;
        RECT  11.810 3.285 12.070 3.940 ;
        RECT  11.080 3.440 11.810 3.940 ;
        RECT  10.820 3.285 11.080 3.940 ;
        RECT  10.280 3.440 10.820 3.940 ;
        RECT  10.020 3.285 10.280 3.940 ;
        RECT  9.370 3.440 10.020 3.940 ;
        RECT  9.110 3.285 9.370 3.940 ;
        RECT  8.305 3.440 9.110 3.940 ;
        RECT  8.045 3.285 8.305 3.940 ;
        RECT  1.735 3.440 8.045 3.940 ;
        RECT  1.475 3.285 1.735 3.940 ;
        RECT  0.785 3.440 1.475 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.840 1.475 15.940 1.735 ;
        RECT  15.680 0.690 15.840 1.735 ;
        RECT  14.780 0.690 15.680 0.850 ;
        RECT  15.190 1.035 15.290 1.295 ;
        RECT  15.190 1.955 15.290 2.555 ;
        RECT  15.030 1.035 15.190 2.555 ;
        RECT  14.805 1.475 15.030 1.735 ;
        RECT  14.625 0.590 14.780 1.215 ;
        RECT  14.465 0.590 14.625 2.990 ;
        RECT  13.730 0.590 14.465 0.750 ;
        RECT  14.365 2.050 14.465 2.990 ;
        RECT  14.115 0.955 14.240 1.215 ;
        RECT  13.955 0.955 14.115 3.105 ;
        RECT  13.855 2.055 13.955 3.105 ;
        RECT  10.750 2.945 13.855 3.105 ;
        RECT  13.630 0.590 13.730 1.210 ;
        RECT  13.470 0.590 13.630 2.765 ;
        RECT  13.345 2.165 13.470 2.765 ;
        RECT  12.585 2.605 13.345 2.765 ;
        RECT  13.120 0.585 13.220 1.210 ;
        RECT  12.960 0.585 13.120 2.425 ;
        RECT  11.840 0.585 12.960 0.745 ;
        RECT  12.835 2.165 12.960 2.425 ;
        RECT  12.585 0.955 12.710 1.215 ;
        RECT  12.425 0.955 12.585 2.765 ;
        RECT  12.325 2.165 12.425 2.765 ;
        RECT  11.680 0.585 11.840 2.325 ;
        RECT  11.540 0.935 11.680 1.195 ;
        RECT  11.670 2.165 11.680 2.325 ;
        RECT  11.410 2.165 11.670 2.765 ;
        RECT  11.240 1.645 11.500 1.905 ;
        RECT  11.195 1.645 11.240 1.805 ;
        RECT  11.035 0.585 11.195 1.805 ;
        RECT  6.850 0.585 11.035 0.745 ;
        RECT  10.750 1.035 10.850 1.295 ;
        RECT  10.590 1.035 10.750 3.105 ;
        RECT  10.420 2.315 10.590 2.915 ;
        RECT  10.155 1.595 10.380 1.855 ;
        RECT  10.120 1.595 10.155 3.105 ;
        RECT  9.995 1.695 10.120 3.105 ;
        RECT  7.695 2.945 9.995 3.105 ;
        RECT  9.670 0.925 9.910 1.185 ;
        RECT  9.670 2.165 9.770 2.765 ;
        RECT  9.650 0.925 9.670 2.765 ;
        RECT  9.510 0.975 9.650 2.765 ;
        RECT  8.820 0.975 9.510 1.135 ;
        RECT  8.820 2.605 9.510 2.765 ;
        RECT  8.560 0.925 8.820 1.185 ;
        RECT  8.560 2.170 8.820 2.765 ;
        RECT  7.355 2.605 8.560 2.765 ;
        RECT  7.700 1.035 7.870 1.295 ;
        RECT  7.700 2.105 7.755 2.365 ;
        RECT  7.540 1.035 7.700 2.365 ;
        RECT  7.535 2.945 7.695 3.220 ;
        RECT  7.405 1.500 7.540 1.760 ;
        RECT  7.495 2.105 7.540 2.365 ;
        RECT  3.395 3.060 7.535 3.220 ;
        RECT  7.190 1.020 7.360 1.280 ;
        RECT  7.255 2.605 7.355 2.880 ;
        RECT  7.190 1.940 7.255 2.880 ;
        RECT  7.095 1.020 7.190 2.880 ;
        RECT  7.030 1.020 7.095 2.100 ;
        RECT  5.255 2.720 7.095 2.880 ;
        RECT  6.745 0.585 6.850 1.280 ;
        RECT  6.745 2.280 6.845 2.540 ;
        RECT  6.690 0.585 6.745 2.540 ;
        RECT  6.585 1.020 6.690 2.540 ;
        RECT  5.765 2.380 6.585 2.540 ;
        RECT  6.205 0.920 6.340 1.180 ;
        RECT  6.205 2.040 6.305 2.200 ;
        RECT  6.045 0.650 6.205 2.200 ;
        RECT  4.890 0.650 6.045 0.810 ;
        RECT  5.730 0.995 5.830 1.255 ;
        RECT  5.730 2.280 5.765 2.540 ;
        RECT  5.570 0.995 5.730 2.540 ;
        RECT  5.505 2.280 5.570 2.540 ;
        RECT  5.205 1.195 5.290 1.455 ;
        RECT  5.205 2.620 5.255 2.880 ;
        RECT  5.045 1.195 5.205 2.880 ;
        RECT  5.030 1.195 5.045 1.455 ;
        RECT  4.995 2.620 5.045 2.880 ;
        RECT  3.835 2.720 4.995 2.880 ;
        RECT  4.790 0.650 4.890 0.945 ;
        RECT  4.790 2.115 4.855 2.375 ;
        RECT  4.630 0.470 4.790 2.375 ;
        RECT  2.715 0.470 4.630 0.630 ;
        RECT  4.595 2.115 4.630 2.375 ;
        RECT  4.280 0.810 4.380 1.070 ;
        RECT  4.280 2.255 4.345 2.515 ;
        RECT  4.120 0.810 4.280 2.515 ;
        RECT  3.395 0.810 4.120 0.970 ;
        RECT  4.085 2.255 4.120 2.515 ;
        RECT  3.735 1.150 3.835 1.310 ;
        RECT  3.735 2.620 3.835 2.880 ;
        RECT  3.575 1.150 3.735 2.880 ;
        RECT  3.235 0.810 3.395 3.220 ;
        RECT  3.015 0.810 3.235 1.070 ;
        RECT  2.845 2.715 3.235 2.975 ;
        RECT  2.555 0.470 2.715 2.145 ;
        RECT  2.455 0.470 2.555 1.095 ;
        RECT  2.285 1.985 2.555 2.145 ;
        RECT  1.335 0.935 2.455 1.095 ;
        RECT  2.215 1.275 2.375 1.805 ;
        RECT  2.025 1.985 2.285 2.330 ;
        RECT  0.385 1.275 2.215 1.435 ;
        RECT  1.335 2.170 2.025 2.330 ;
        RECT  1.075 0.495 1.335 1.095 ;
        RECT  1.075 2.170 1.335 2.430 ;
        RECT  0.285 0.855 0.385 1.435 ;
        RECT  0.285 2.055 0.385 2.315 ;
        RECT  0.125 0.855 0.285 2.315 ;
    END
END BMXX4

MACRO BMXX2
    CLASS CORE ;
    FOREIGN BMXX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.525 2.555 9.805 3.230 ;
        RECT  9.325 2.930 9.525 3.220 ;
        END
        ANTENNAGATEAREA     0.2951 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 1.290 6.775 1.785 ;
        RECT  6.475 1.440 6.565 1.785 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.905 0.695 10.915 0.945 ;
        RECT  10.905 2.110 10.915 2.585 ;
        RECT  10.745 0.695 10.905 2.915 ;
        RECT  10.730 0.695 10.745 1.355 ;
        RECT  10.730 1.925 10.745 2.915 ;
        RECT  10.645 0.695 10.730 1.295 ;
        RECT  10.645 1.975 10.730 2.915 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.645 1.290 5.855 1.815 ;
        RECT  5.435 1.555 5.645 1.815 ;
        END
        ANTENNAGATEAREA     0.2275 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.455 1.490 2.615 2.780 ;
        RECT  2.105 2.620 2.455 2.780 ;
        RECT  2.005 2.620 2.105 2.880 ;
        RECT  1.845 2.620 2.005 3.105 ;
        RECT  0.795 2.945 1.845 3.105 ;
        RECT  0.585 1.615 0.795 3.105 ;
        RECT  0.475 1.615 0.585 1.875 ;
        END
        ANTENNAGATEAREA     0.2275 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.975 1.615 1.410 1.990 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.345 -0.250 11.040 0.250 ;
        RECT  10.085 -0.250 10.345 0.405 ;
        RECT  7.845 -0.250 10.085 0.250 ;
        RECT  7.585 -0.250 7.845 0.405 ;
        RECT  6.795 -0.250 7.585 0.250 ;
        RECT  5.735 -0.250 6.795 0.405 ;
        RECT  1.765 -0.250 5.735 0.250 ;
        RECT  1.505 -0.250 1.765 0.405 ;
        RECT  0.815 -0.250 1.505 0.250 ;
        RECT  0.555 -0.250 0.815 0.800 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.395 3.440 11.040 3.940 ;
        RECT  10.135 2.275 10.395 3.940 ;
        RECT  7.705 3.440 10.135 3.940 ;
        RECT  7.445 3.285 7.705 3.940 ;
        RECT  6.795 3.440 7.445 3.940 ;
        RECT  5.735 3.285 6.795 3.940 ;
        RECT  5.355 3.440 5.735 3.940 ;
        RECT  3.395 3.390 5.355 3.940 ;
        RECT  1.735 3.440 3.395 3.940 ;
        RECT  1.475 3.285 1.735 3.940 ;
        RECT  0.785 3.440 1.475 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.465 1.475 10.545 1.735 ;
        RECT  10.305 0.685 10.465 1.735 ;
        RECT  8.895 0.685 10.305 0.845 ;
        RECT  9.865 1.035 9.915 1.295 ;
        RECT  9.705 1.035 9.865 2.355 ;
        RECT  9.655 1.035 9.705 1.295 ;
        RECT  9.595 1.725 9.705 2.355 ;
        RECT  9.455 1.725 9.595 1.985 ;
        RECT  9.275 1.035 9.405 1.295 ;
        RECT  9.145 1.035 9.275 2.555 ;
        RECT  9.115 1.035 9.145 2.905 ;
        RECT  8.985 1.955 9.115 2.905 ;
        RECT  7.305 2.745 8.985 2.905 ;
        RECT  8.765 0.685 8.895 1.285 ;
        RECT  8.635 0.685 8.765 2.555 ;
        RECT  8.605 1.125 8.635 2.555 ;
        RECT  8.505 1.955 8.605 2.555 ;
        RECT  8.255 0.695 8.385 1.295 ;
        RECT  8.125 0.695 8.255 2.555 ;
        RECT  8.095 1.135 8.125 2.555 ;
        RECT  7.995 1.955 8.095 2.555 ;
        RECT  7.745 0.655 7.905 1.665 ;
        RECT  4.485 0.655 7.745 0.815 ;
        RECT  7.395 1.135 7.555 2.465 ;
        RECT  7.305 1.135 7.395 1.295 ;
        RECT  7.305 2.305 7.395 2.465 ;
        RECT  7.045 1.035 7.305 1.295 ;
        RECT  7.045 2.305 7.305 2.905 ;
        RECT  7.115 1.475 7.215 1.735 ;
        RECT  6.955 1.475 7.115 2.125 ;
        RECT  6.735 1.965 6.955 2.125 ;
        RECT  6.575 1.965 6.735 2.995 ;
        RECT  5.385 2.835 6.575 2.995 ;
        RECT  6.295 2.055 6.395 2.655 ;
        RECT  6.295 1.000 6.345 1.260 ;
        RECT  6.135 1.000 6.295 2.655 ;
        RECT  5.045 2.495 6.135 2.655 ;
        RECT  5.185 1.995 5.445 2.255 ;
        RECT  5.165 1.035 5.385 1.295 ;
        RECT  5.225 2.835 5.385 3.105 ;
        RECT  2.955 2.945 5.225 3.105 ;
        RECT  5.165 1.995 5.185 2.155 ;
        RECT  5.005 1.035 5.165 2.155 ;
        RECT  4.825 2.495 5.045 2.765 ;
        RECT  4.665 1.035 4.825 2.765 ;
        RECT  3.625 2.605 4.665 2.765 ;
        RECT  4.325 0.655 4.485 2.425 ;
        RECT  4.075 1.035 4.325 1.295 ;
        RECT  3.775 1.955 4.025 2.215 ;
        RECT  3.775 1.035 3.825 1.295 ;
        RECT  3.765 1.035 3.775 2.215 ;
        RECT  3.725 1.035 3.765 2.165 ;
        RECT  3.615 0.470 3.725 2.165 ;
        RECT  3.365 2.505 3.625 2.765 ;
        RECT  3.565 0.470 3.615 1.295 ;
        RECT  2.290 0.470 3.565 0.630 ;
        RECT  3.320 2.505 3.365 2.665 ;
        RECT  3.160 0.810 3.320 2.665 ;
        RECT  3.055 0.810 3.160 0.970 ;
        RECT  2.805 1.150 2.955 3.105 ;
        RECT  2.795 0.960 2.805 3.105 ;
        RECT  2.545 0.960 2.795 1.310 ;
        RECT  2.275 0.470 2.290 1.070 ;
        RECT  2.245 0.470 2.275 2.330 ;
        RECT  2.130 0.470 2.245 2.440 ;
        RECT  2.115 0.810 2.130 2.440 ;
        RECT  2.030 0.810 2.115 1.095 ;
        RECT  1.985 2.170 2.115 2.440 ;
        RECT  1.365 0.935 2.030 1.095 ;
        RECT  1.335 2.170 1.985 2.330 ;
        RECT  1.775 1.275 1.935 1.985 ;
        RECT  0.385 1.275 1.775 1.435 ;
        RECT  1.105 0.835 1.365 1.095 ;
        RECT  1.075 2.170 1.335 2.765 ;
        RECT  0.285 1.035 0.385 1.435 ;
        RECT  0.285 2.095 0.385 2.355 ;
        RECT  0.125 1.035 0.285 2.355 ;
    END
END BMXX2

MACRO BENCX4
    CLASS CORE ;
    FOREIGN BENCX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.745 1.290 23.795 2.085 ;
        RECT  23.585 0.955 23.745 2.085 ;
        RECT  23.465 0.955 23.585 1.215 ;
        RECT  20.225 1.925 23.585 2.085 ;
        RECT  22.645 1.005 23.465 1.165 ;
        RECT  22.385 0.955 22.645 1.215 ;
        RECT  21.565 1.005 22.385 1.165 ;
        RECT  21.305 0.955 21.565 1.215 ;
        RECT  20.485 1.005 21.305 1.165 ;
        RECT  20.225 0.955 20.485 1.215 ;
        END
        ANTENNADIFFAREA     3.1312 ;
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  33.495 0.695 33.755 1.295 ;
        RECT  33.480 1.035 33.495 1.295 ;
        RECT  33.220 1.035 33.480 2.430 ;
        RECT  32.735 1.035 33.220 1.295 ;
        RECT  32.860 2.170 33.220 2.430 ;
        RECT  32.600 2.170 32.860 3.215 ;
        RECT  32.475 0.695 32.735 1.295 ;
        RECT  31.840 2.170 32.600 2.430 ;
        RECT  31.715 1.035 32.475 1.295 ;
        RECT  31.580 2.170 31.840 3.215 ;
        RECT  31.455 0.695 31.715 1.295 ;
        RECT  30.820 2.170 31.580 2.430 ;
        RECT  30.695 1.035 31.455 1.295 ;
        RECT  30.560 2.170 30.820 3.215 ;
        RECT  30.435 0.695 30.695 1.295 ;
        RECT  29.800 2.170 30.560 2.430 ;
        RECT  29.540 2.170 29.800 3.215 ;
        END
        ANTENNADIFFAREA     3.2832 ;
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.170 2.945 24.645 3.105 ;
        RECT  16.945 2.945 17.170 3.215 ;
        RECT  14.285 3.055 16.945 3.215 ;
        RECT  14.125 2.945 14.285 3.215 ;
        RECT  9.125 2.945 14.125 3.105 ;
        RECT  9.075 2.930 9.125 3.190 ;
        RECT  8.865 2.930 9.075 3.220 ;
        END
        ANTENNAGATEAREA     0.4082 ;
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.830 2.590 14.285 2.750 ;
        RECT  8.670 2.170 8.830 2.750 ;
        RECT  7.975 2.170 8.670 2.330 ;
        RECT  7.815 1.760 7.975 2.330 ;
        RECT  7.670 1.760 7.815 2.020 ;
        RECT  6.775 1.810 7.670 1.970 ;
        RECT  6.625 1.700 6.775 1.990 ;
        RECT  6.565 1.700 6.625 2.020 ;
        RECT  6.465 1.760 6.565 2.020 ;
        END
        ANTENNAGATEAREA     1.1648 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.975 1.360 12.235 1.620 ;
        RECT  11.925 1.360 11.975 1.520 ;
        RECT  11.765 0.585 11.925 1.520 ;
        RECT  10.245 0.585 11.765 0.745 ;
        RECT  10.085 0.585 10.245 1.455 ;
        RECT  9.970 1.290 10.085 1.455 ;
        RECT  7.235 1.295 9.970 1.455 ;
        RECT  7.025 1.290 7.235 1.580 ;
        RECT  6.480 1.295 7.025 1.455 ;
        END
        ANTENNAGATEAREA     1.1687 ;
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.955 2.745 4.015 2.995 ;
        RECT  3.695 0.695 3.955 1.295 ;
        RECT  3.695 2.165 3.955 3.105 ;
        RECT  2.935 1.035 3.695 1.295 ;
        RECT  2.935 2.165 3.695 2.425 ;
        RECT  2.675 0.695 2.935 1.295 ;
        RECT  2.675 2.165 2.935 3.105 ;
        RECT  1.915 1.035 2.675 1.295 ;
        RECT  1.915 2.165 2.675 2.425 ;
        RECT  1.655 0.695 1.915 1.295 ;
        RECT  1.655 2.165 1.915 3.105 ;
        RECT  0.895 1.035 1.655 1.295 ;
        RECT  1.075 2.165 1.655 2.425 ;
        RECT  0.895 2.110 1.075 2.425 ;
        RECT  0.635 0.695 0.895 3.180 ;
        RECT  0.585 1.105 0.635 2.995 ;
        END
        ANTENNADIFFAREA     3.2832 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  34.265 -0.250 34.500 0.250 ;
        RECT  34.005 -0.250 34.265 1.290 ;
        RECT  33.245 -0.250 34.005 0.250 ;
        RECT  32.985 -0.250 33.245 0.735 ;
        RECT  32.225 -0.250 32.985 0.250 ;
        RECT  31.965 -0.250 32.225 0.735 ;
        RECT  31.205 -0.250 31.965 0.250 ;
        RECT  30.945 -0.250 31.205 0.735 ;
        RECT  30.185 -0.250 30.945 0.250 ;
        RECT  29.925 -0.250 30.185 1.115 ;
        RECT  29.165 -0.250 29.925 0.250 ;
        RECT  28.905 -0.250 29.165 1.115 ;
        RECT  28.255 -0.250 28.905 0.250 ;
        RECT  27.995 -0.250 28.255 0.405 ;
        RECT  27.165 -0.250 27.995 0.250 ;
        RECT  26.905 -0.250 27.165 0.405 ;
        RECT  26.085 -0.250 26.905 0.250 ;
        RECT  25.825 -0.250 26.085 0.405 ;
        RECT  24.265 -0.250 25.825 0.250 ;
        RECT  24.005 -0.250 24.265 0.405 ;
        RECT  23.185 -0.250 24.005 0.250 ;
        RECT  22.925 -0.250 23.185 0.405 ;
        RECT  22.105 -0.250 22.925 0.250 ;
        RECT  21.845 -0.250 22.105 0.405 ;
        RECT  21.025 -0.250 21.845 0.250 ;
        RECT  20.765 -0.250 21.025 0.405 ;
        RECT  19.945 -0.250 20.765 0.250 ;
        RECT  19.685 -0.250 19.945 0.405 ;
        RECT  19.005 -0.250 19.685 0.250 ;
        RECT  18.745 -0.250 19.005 0.405 ;
        RECT  17.925 -0.250 18.745 0.250 ;
        RECT  17.665 -0.250 17.925 0.405 ;
        RECT  15.055 -0.250 17.665 0.250 ;
        RECT  14.795 -0.250 15.055 0.405 ;
        RECT  13.955 -0.250 14.795 0.250 ;
        RECT  13.695 -0.250 13.955 0.405 ;
        RECT  13.045 -0.250 13.695 0.250 ;
        RECT  12.785 -0.250 13.045 1.145 ;
        RECT  11.985 -0.250 12.785 0.250 ;
        RECT  11.725 -0.250 11.985 0.405 ;
        RECT  11.035 -0.250 11.725 0.250 ;
        RECT  10.775 -0.250 11.035 0.405 ;
        RECT  8.535 -0.250 10.775 0.250 ;
        RECT  8.275 -0.250 8.535 0.405 ;
        RECT  7.450 -0.250 8.275 0.250 ;
        RECT  7.190 -0.250 7.450 0.405 ;
        RECT  6.400 -0.250 7.190 0.250 ;
        RECT  6.140 -0.250 6.400 0.755 ;
        RECT  5.485 -0.250 6.140 0.250 ;
        RECT  5.225 -0.250 5.485 0.875 ;
        RECT  4.465 -0.250 5.225 0.250 ;
        RECT  4.205 -0.250 4.465 0.880 ;
        RECT  3.445 -0.250 4.205 0.250 ;
        RECT  3.185 -0.250 3.445 0.785 ;
        RECT  2.425 -0.250 3.185 0.250 ;
        RECT  2.165 -0.250 2.425 0.735 ;
        RECT  1.405 -0.250 2.165 0.250 ;
        RECT  1.145 -0.250 1.405 0.735 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.075 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  33.370 3.440 34.500 3.940 ;
        RECT  33.110 2.615 33.370 3.940 ;
        RECT  32.350 3.440 33.110 3.940 ;
        RECT  32.090 2.615 32.350 3.940 ;
        RECT  31.330 3.440 32.090 3.940 ;
        RECT  31.070 2.615 31.330 3.940 ;
        RECT  30.310 3.440 31.070 3.940 ;
        RECT  30.050 2.615 30.310 3.940 ;
        RECT  29.290 3.440 30.050 3.940 ;
        RECT  29.030 2.465 29.290 3.940 ;
        RECT  28.270 3.440 29.030 3.940 ;
        RECT  28.010 2.465 28.270 3.940 ;
        RECT  27.250 3.440 28.010 3.940 ;
        RECT  26.990 2.255 27.250 3.940 ;
        RECT  25.575 3.440 26.990 3.940 ;
        RECT  25.315 3.285 25.575 3.940 ;
        RECT  24.275 3.440 25.315 3.940 ;
        RECT  24.015 3.285 24.275 3.940 ;
        RECT  23.185 3.440 24.015 3.940 ;
        RECT  22.925 3.285 23.185 3.940 ;
        RECT  22.105 3.440 22.925 3.940 ;
        RECT  21.845 3.285 22.105 3.940 ;
        RECT  21.025 3.440 21.845 3.940 ;
        RECT  20.765 3.285 21.025 3.940 ;
        RECT  19.945 3.440 20.765 3.940 ;
        RECT  19.685 3.285 19.945 3.940 ;
        RECT  19.015 3.440 19.685 3.940 ;
        RECT  18.755 3.285 19.015 3.940 ;
        RECT  17.840 3.440 18.755 3.940 ;
        RECT  17.580 3.285 17.840 3.940 ;
        RECT  13.915 3.440 17.580 3.940 ;
        RECT  13.655 3.285 13.915 3.940 ;
        RECT  13.115 3.440 13.655 3.940 ;
        RECT  12.855 3.285 13.115 3.940 ;
        RECT  12.015 3.440 12.855 3.940 ;
        RECT  11.755 3.285 12.015 3.940 ;
        RECT  10.570 3.440 11.755 3.940 ;
        RECT  10.310 3.285 10.570 3.940 ;
        RECT  9.770 3.440 10.310 3.940 ;
        RECT  9.510 3.285 9.770 3.940 ;
        RECT  8.145 3.440 9.510 3.940 ;
        RECT  7.885 2.850 8.145 3.940 ;
        RECT  6.505 3.440 7.885 3.940 ;
        RECT  6.245 2.540 6.505 3.940 ;
        RECT  5.485 3.440 6.245 3.940 ;
        RECT  5.225 2.415 5.485 3.940 ;
        RECT  4.465 3.440 5.225 3.940 ;
        RECT  4.205 2.415 4.465 3.940 ;
        RECT  3.445 3.440 4.205 3.940 ;
        RECT  3.185 2.615 3.445 3.940 ;
        RECT  2.425 3.440 3.185 3.940 ;
        RECT  2.165 2.615 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.615 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  30.025 1.585 33.005 1.845 ;
        RECT  29.675 1.635 30.025 1.795 ;
        RECT  29.415 0.595 29.675 1.795 ;
        RECT  29.375 0.815 29.415 1.795 ;
        RECT  28.685 1.635 29.375 1.795 ;
        RECT  28.685 2.125 28.780 3.065 ;
        RECT  28.525 0.935 28.685 3.065 ;
        RECT  28.395 0.935 28.525 1.195 ;
        RECT  28.520 2.125 28.525 3.065 ;
        RECT  27.760 2.125 28.520 2.285 ;
        RECT  28.045 1.635 28.340 1.900 ;
        RECT  27.885 0.620 28.045 1.900 ;
        RECT  24.915 0.620 27.885 0.780 ;
        RECT  27.740 1.635 27.885 1.900 ;
        RECT  27.500 2.125 27.760 3.065 ;
        RECT  26.595 1.740 27.740 1.900 ;
        RECT  24.665 0.960 27.705 1.120 ;
        RECT  27.125 1.300 27.385 1.560 ;
        RECT  25.985 1.365 27.125 1.525 ;
        RECT  26.435 1.740 26.595 2.410 ;
        RECT  26.425 2.250 26.435 2.410 ;
        RECT  26.165 2.250 26.425 3.190 ;
        RECT  25.985 1.810 26.255 2.070 ;
        RECT  24.985 2.665 26.165 2.825 ;
        RECT  25.825 1.365 25.985 2.485 ;
        RECT  24.175 1.365 25.825 1.525 ;
        RECT  24.475 2.325 25.825 2.485 ;
        RECT  25.475 1.840 25.635 2.100 ;
        RECT  24.135 1.890 25.475 2.050 ;
        RECT  24.825 2.665 24.985 2.925 ;
        RECT  24.405 0.925 24.665 1.185 ;
        RECT  24.315 2.325 24.475 2.765 ;
        RECT  16.765 2.605 24.315 2.765 ;
        RECT  24.015 0.585 24.175 1.525 ;
        RECT  23.975 1.890 24.135 2.425 ;
        RECT  13.555 0.585 24.015 0.745 ;
        RECT  16.765 2.265 23.975 2.425 ;
        RECT  19.555 1.465 23.295 1.725 ;
        RECT  19.545 1.465 19.555 2.085 ;
        RECT  19.395 0.955 19.545 2.085 ;
        RECT  19.385 0.955 19.395 1.675 ;
        RECT  18.215 1.925 19.395 2.085 ;
        RECT  19.285 0.955 19.385 1.215 ;
        RECT  18.465 1.055 19.285 1.215 ;
        RECT  17.895 1.485 18.975 1.745 ;
        RECT  18.205 0.955 18.465 1.215 ;
        RECT  17.735 0.925 17.895 2.085 ;
        RECT  15.705 0.925 17.735 1.085 ;
        RECT  16.255 1.925 17.735 2.085 ;
        RECT  15.805 1.265 17.555 1.425 ;
        RECT  16.505 2.605 16.765 2.875 ;
        RECT  14.465 2.715 16.505 2.875 ;
        RECT  16.095 1.925 16.255 2.530 ;
        RECT  14.975 2.370 16.095 2.530 ;
        RECT  15.645 1.265 15.805 2.190 ;
        RECT  15.470 1.265 15.645 1.425 ;
        RECT  14.520 2.030 15.645 2.190 ;
        RECT  15.310 0.955 15.470 1.425 ;
        RECT  14.035 1.660 15.465 1.820 ;
        RECT  14.245 0.955 15.310 1.115 ;
        RECT  14.360 2.030 14.520 2.410 ;
        RECT  13.255 2.250 14.360 2.410 ;
        RECT  13.875 1.660 14.035 2.070 ;
        RECT  12.915 1.910 13.875 2.070 ;
        RECT  13.555 1.470 13.695 1.730 ;
        RECT  13.395 0.585 13.555 1.730 ;
        RECT  13.295 0.935 13.395 1.730 ;
        RECT  12.575 1.520 13.295 1.730 ;
        RECT  12.755 1.910 12.915 2.410 ;
        RECT  10.925 2.250 12.755 2.410 ;
        RECT  12.415 0.580 12.575 2.070 ;
        RECT  12.275 0.580 12.415 1.180 ;
        RECT  11.355 1.910 12.415 2.070 ;
        RECT  11.325 0.925 11.585 1.185 ;
        RECT  10.925 1.025 11.325 1.185 ;
        RECT  10.765 1.025 10.925 2.410 ;
        RECT  9.910 2.250 10.765 2.410 ;
        RECT  10.425 0.925 10.585 2.070 ;
        RECT  9.170 1.910 10.425 2.070 ;
        RECT  9.745 0.795 9.905 1.095 ;
        RECT  6.285 0.935 9.745 1.095 ;
        RECT  7.995 0.595 9.445 0.755 ;
        RECT  9.010 1.830 9.170 2.215 ;
        RECT  8.485 1.830 9.010 1.990 ;
        RECT  8.485 2.940 8.685 3.100 ;
        RECT  8.225 1.730 8.485 1.990 ;
        RECT  8.325 2.510 8.485 3.100 ;
        RECT  7.325 2.510 8.325 2.670 ;
        RECT  7.735 0.495 7.995 0.755 ;
        RECT  6.910 0.595 7.735 0.755 ;
        RECT  7.065 2.150 7.325 3.090 ;
        RECT  6.285 2.200 7.065 2.360 ;
        RECT  6.650 0.495 6.910 0.755 ;
        RECT  6.125 0.935 6.285 2.360 ;
        RECT  5.490 1.545 6.125 1.705 ;
        RECT  5.785 1.035 5.945 1.295 ;
        RECT  5.785 1.955 5.945 2.895 ;
        RECT  4.975 1.135 5.785 1.295 ;
        RECT  4.975 2.075 5.785 2.235 ;
        RECT  4.550 1.495 5.490 1.755 ;
        RECT  4.715 0.695 4.975 1.295 ;
        RECT  4.715 2.075 4.975 3.015 ;
        RECT  4.295 1.135 4.715 1.295 ;
        RECT  4.295 2.075 4.715 2.235 ;
        RECT  4.135 1.135 4.295 2.235 ;
        RECT  1.155 1.475 4.135 1.735 ;
    END
END BENCX4

MACRO BENCX2
    CLASS CORE ;
    FOREIGN BENCX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.320 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.755 1.920 13.425 2.080 ;
        RECT  13.090 0.935 13.350 1.195 ;
        RECT  12.335 0.985 13.090 1.145 ;
        RECT  12.545 1.700 12.755 2.080 ;
        RECT  12.335 1.920 12.545 2.080 ;
        RECT  12.270 0.985 12.335 2.080 ;
        RECT  12.175 0.935 12.270 2.080 ;
        RECT  12.010 0.935 12.175 1.195 ;
        RECT  12.085 1.920 12.175 2.080 ;
        END
        ANTENNADIFFAREA     1.5504 ;
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.985 1.700 19.195 1.990 ;
        RECT  18.735 1.765 18.985 1.925 ;
        RECT  18.700 1.100 18.735 2.585 ;
        RECT  18.685 0.915 18.700 2.585 ;
        RECT  18.525 0.695 18.685 2.930 ;
        RECT  18.425 0.695 18.525 1.420 ;
        RECT  18.425 1.990 18.525 2.930 ;
        RECT  17.665 1.260 18.425 1.420 ;
        RECT  17.665 1.990 18.425 2.150 ;
        RECT  17.405 0.695 17.665 1.420 ;
        RECT  17.405 1.990 17.665 2.930 ;
        END
        ANTENNADIFFAREA     1.6546 ;
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.305 2.930 15.515 3.220 ;
        RECT  11.005 2.945 15.305 3.105 ;
        RECT  10.845 2.945 11.005 3.220 ;
        RECT  8.525 3.060 10.845 3.220 ;
        RECT  8.365 2.945 8.525 3.220 ;
        RECT  6.285 2.945 8.365 3.105 ;
        END
        ANTENNAGATEAREA     0.2041 ;
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 1.975 8.585 2.135 ;
        RECT  7.870 1.975 8.030 2.765 ;
        RECT  6.015 2.605 7.870 2.765 ;
        RECT  5.855 2.605 6.015 3.205 ;
        RECT  4.475 2.605 5.855 2.765 ;
        RECT  4.315 1.680 4.475 2.765 ;
        RECT  4.265 1.680 4.315 2.400 ;
        RECT  4.155 1.680 4.265 1.840 ;
        END
        ANTENNAGATEAREA     0.5863 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 0.505 6.955 0.665 ;
        RECT  6.155 0.505 6.315 0.970 ;
        RECT  6.130 0.695 6.155 0.970 ;
        RECT  5.235 0.810 6.130 0.970 ;
        RECT  5.075 0.810 5.235 1.430 ;
        RECT  3.850 1.270 5.075 1.430 ;
        RECT  3.590 1.270 3.850 1.820 ;
        RECT  3.345 1.270 3.590 1.580 ;
        END
        ANTENNAGATEAREA     0.5850 ;
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 0.695 1.915 1.415 ;
        RECT  1.655 2.125 1.915 3.065 ;
        RECT  0.895 1.255 1.655 1.415 ;
        RECT  1.070 2.125 1.655 2.285 ;
        RECT  0.895 2.125 1.070 2.400 ;
        RECT  0.795 0.695 0.895 1.415 ;
        RECT  0.795 2.125 0.895 3.065 ;
        RECT  0.635 0.695 0.795 3.065 ;
        RECT  0.585 1.105 0.635 2.590 ;
        END
        ANTENNADIFFAREA     1.6416 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.195 -0.250 19.320 0.250 ;
        RECT  18.935 -0.250 19.195 1.075 ;
        RECT  18.175 -0.250 18.935 0.250 ;
        RECT  17.915 -0.250 18.175 1.075 ;
        RECT  17.065 -0.250 17.915 0.250 ;
        RECT  16.805 -0.250 17.065 0.405 ;
        RECT  16.290 -0.250 16.805 0.250 ;
        RECT  16.030 -0.250 16.290 0.405 ;
        RECT  15.200 -0.250 16.030 0.250 ;
        RECT  14.940 -0.250 15.200 0.405 ;
        RECT  13.890 -0.250 14.940 0.250 ;
        RECT  13.630 -0.250 13.890 0.405 ;
        RECT  12.810 -0.250 13.630 0.250 ;
        RECT  12.550 -0.250 12.810 0.405 ;
        RECT  11.730 -0.250 12.550 0.250 ;
        RECT  11.470 -0.250 11.730 0.405 ;
        RECT  10.650 -0.250 11.470 0.250 ;
        RECT  10.390 -0.250 10.650 0.405 ;
        RECT  8.400 -0.250 10.390 0.250 ;
        RECT  8.140 -0.250 8.400 0.405 ;
        RECT  7.300 -0.250 8.140 0.250 ;
        RECT  7.140 -0.250 7.300 0.755 ;
        RECT  5.945 -0.250 7.140 0.250 ;
        RECT  5.685 -0.250 5.945 0.405 ;
        RECT  4.495 -0.250 5.685 0.250 ;
        RECT  4.235 -0.250 4.495 0.405 ;
        RECT  3.445 -0.250 4.235 0.250 ;
        RECT  3.185 -0.250 3.445 0.735 ;
        RECT  2.425 -0.250 3.185 0.250 ;
        RECT  2.165 -0.250 2.425 0.830 ;
        RECT  1.405 -0.250 2.165 0.250 ;
        RECT  1.145 -0.250 1.405 1.075 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.075 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.195 3.440 19.320 3.940 ;
        RECT  18.935 2.265 19.195 3.940 ;
        RECT  18.175 3.440 18.935 3.940 ;
        RECT  17.915 2.435 18.175 3.940 ;
        RECT  17.055 3.440 17.915 3.940 ;
        RECT  16.795 3.285 17.055 3.940 ;
        RECT  16.155 3.440 16.795 3.940 ;
        RECT  15.895 2.800 16.155 3.940 ;
        RECT  15.045 3.440 15.895 3.940 ;
        RECT  14.785 3.285 15.045 3.940 ;
        RECT  13.965 3.440 14.785 3.940 ;
        RECT  13.705 3.285 13.965 3.940 ;
        RECT  12.885 3.440 13.705 3.940 ;
        RECT  12.625 3.285 12.885 3.940 ;
        RECT  11.795 3.440 12.625 3.940 ;
        RECT  11.535 3.285 11.795 3.940 ;
        RECT  7.775 3.440 11.535 3.940 ;
        RECT  7.515 3.285 7.775 3.940 ;
        RECT  6.915 3.440 7.515 3.940 ;
        RECT  6.655 3.285 6.915 3.940 ;
        RECT  5.645 3.440 6.655 3.940 ;
        RECT  5.485 2.945 5.645 3.940 ;
        RECT  4.585 3.440 5.485 3.940 ;
        RECT  4.325 3.285 4.585 3.940 ;
        RECT  3.485 3.440 4.325 3.940 ;
        RECT  3.225 3.285 3.485 3.940 ;
        RECT  2.425 3.440 3.225 3.940 ;
        RECT  2.165 2.615 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.610 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.795 1.605 18.165 1.765 ;
        RECT  16.695 0.940 16.795 2.120 ;
        RECT  16.635 0.940 16.695 2.560 ;
        RECT  16.435 0.940 16.635 1.200 ;
        RECT  16.435 1.960 16.635 2.560 ;
        RECT  16.185 1.405 16.445 1.665 ;
        RECT  15.875 1.455 16.185 1.615 ;
        RECT  15.755 0.925 15.875 2.445 ;
        RECT  15.715 0.925 15.755 2.545 ;
        RECT  14.290 0.585 15.740 0.745 ;
        RECT  14.540 0.925 15.715 1.085 ;
        RECT  15.495 2.285 15.715 2.545 ;
        RECT  15.375 1.265 15.535 2.105 ;
        RECT  14.445 2.285 15.495 2.445 ;
        RECT  13.740 1.265 15.375 1.425 ;
        RECT  14.105 1.945 15.375 2.105 ;
        RECT  13.765 1.605 15.105 1.765 ;
        RECT  14.285 2.285 14.445 2.545 ;
        RECT  14.130 0.585 14.290 1.085 ;
        RECT  14.030 0.825 14.130 1.085 ;
        RECT  13.945 1.945 14.105 2.765 ;
        RECT  10.665 2.605 13.945 2.765 ;
        RECT  13.605 1.605 13.765 2.420 ;
        RECT  13.580 0.585 13.740 1.425 ;
        RECT  10.665 2.260 13.605 2.420 ;
        RECT  7.865 0.585 13.580 0.745 ;
        RECT  11.835 1.405 11.995 1.665 ;
        RECT  11.400 1.455 11.835 1.615 ;
        RECT  11.350 1.455 11.400 2.075 ;
        RECT  11.240 0.985 11.350 2.075 ;
        RECT  11.190 0.985 11.240 1.615 ;
        RECT  11.135 1.915 11.240 2.075 ;
        RECT  10.930 0.935 11.190 1.195 ;
        RECT  10.505 1.755 10.665 2.420 ;
        RECT  10.505 2.605 10.665 2.880 ;
        RECT  8.705 2.720 10.505 2.880 ;
        RECT  10.325 0.925 10.330 1.085 ;
        RECT  10.165 0.925 10.325 2.540 ;
        RECT  9.190 0.925 10.165 1.085 ;
        RECT  9.215 2.380 10.165 2.540 ;
        RECT  9.825 1.295 9.985 2.200 ;
        RECT  8.975 1.295 9.825 1.455 ;
        RECT  8.995 2.040 9.825 2.200 ;
        RECT  7.685 1.635 9.620 1.795 ;
        RECT  8.835 2.040 8.995 2.475 ;
        RECT  8.815 0.925 8.975 1.455 ;
        RECT  8.370 2.315 8.835 2.475 ;
        RECT  8.680 0.925 8.815 1.085 ;
        RECT  7.865 1.295 8.600 1.455 ;
        RECT  8.210 2.315 8.370 2.765 ;
        RECT  7.705 0.585 7.865 1.455 ;
        RECT  7.700 0.735 7.705 1.455 ;
        RECT  7.600 0.735 7.700 0.995 ;
        RECT  7.345 1.295 7.700 1.455 ;
        RECT  7.525 1.635 7.685 2.425 ;
        RECT  6.680 2.265 7.525 2.425 ;
        RECT  7.185 1.295 7.345 2.085 ;
        RECT  7.085 1.925 7.185 2.085 ;
        RECT  6.680 0.955 6.780 1.215 ;
        RECT  6.520 0.955 6.680 2.425 ;
        RECT  5.975 2.165 6.520 2.425 ;
        RECT  5.575 1.155 5.805 1.315 ;
        RECT  5.415 1.155 5.575 1.775 ;
        RECT  4.835 0.470 5.435 0.630 ;
        RECT  5.085 1.615 5.415 1.775 ;
        RECT  5.085 2.095 5.155 2.355 ;
        RECT  3.705 2.945 5.125 3.105 ;
        RECT  4.925 1.615 5.085 2.355 ;
        RECT  4.695 1.615 4.925 1.875 ;
        RECT  4.895 2.095 4.925 2.355 ;
        RECT  3.105 0.930 4.895 1.090 ;
        RECT  4.675 0.470 4.835 0.745 ;
        RECT  3.695 0.585 4.675 0.745 ;
        RECT  3.705 2.000 3.735 2.600 ;
        RECT  3.545 2.000 3.705 3.105 ;
        RECT  3.475 2.000 3.545 2.600 ;
        RECT  3.410 2.000 3.475 2.160 ;
        RECT  3.250 1.760 3.410 2.160 ;
        RECT  3.105 1.760 3.250 1.920 ;
        RECT  2.945 0.930 3.105 1.920 ;
        RECT  2.695 1.580 2.945 1.740 ;
        RECT  2.765 0.480 2.935 0.740 ;
        RECT  2.885 2.875 2.935 3.135 ;
        RECT  2.725 2.105 2.885 3.135 ;
        RECT  2.605 0.480 2.765 1.175 ;
        RECT  2.255 2.105 2.725 2.265 ;
        RECT  2.675 2.875 2.725 3.135 ;
        RECT  2.435 1.530 2.695 1.790 ;
        RECT  2.255 1.015 2.605 1.175 ;
        RECT  2.095 1.015 2.255 2.265 ;
        RECT  0.985 1.635 2.095 1.795 ;
    END
END BENCX2

MACRO BENCX1
    CLASS CORE ;
    FOREIGN BENCX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.950 0.925 10.110 2.085 ;
        RECT  9.680 0.925 9.950 1.180 ;
        RECT  9.810 1.700 9.950 2.085 ;
        RECT  9.785 1.700 9.810 1.990 ;
        END
        ANTENNADIFFAREA     0.7638 ;
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.085 1.515 14.135 1.990 ;
        RECT  14.000 1.275 14.085 2.190 ;
        RECT  13.925 0.695 14.000 2.970 ;
        RECT  13.740 0.695 13.925 1.435 ;
        RECT  13.740 2.030 13.925 2.970 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.165 2.895 11.375 3.220 ;
        RECT  11.115 2.895 11.165 3.155 ;
        RECT  9.095 2.945 11.115 3.105 ;
        RECT  8.935 2.945 9.095 3.220 ;
        RECT  6.645 3.060 8.935 3.220 ;
        RECT  6.485 2.945 6.645 3.220 ;
        RECT  4.810 2.945 6.485 3.105 ;
        END
        ANTENNAGATEAREA     0.1274 ;
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.865 2.605 6.645 2.765 ;
        RECT  2.865 1.815 2.970 1.975 ;
        RECT  2.705 1.815 2.865 2.765 ;
        RECT  2.425 2.110 2.705 2.400 ;
        END
        ANTENNAGATEAREA     0.2964 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.125 0.585 5.635 0.745 ;
        RECT  3.965 0.585 4.125 1.595 ;
        RECT  2.525 1.435 3.965 1.595 ;
        RECT  2.365 1.435 2.525 1.785 ;
        RECT  2.175 1.525 2.365 1.785 ;
        RECT  2.155 1.525 2.175 1.990 ;
        RECT  1.990 1.575 2.155 1.990 ;
        RECT  1.965 1.700 1.990 1.990 ;
        END
        ANTENNAGATEAREA     0.2951 ;
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.635 0.695 0.895 1.435 ;
        RECT  0.635 1.975 0.895 2.915 ;
        RECT  0.585 1.105 0.635 1.435 ;
        RECT  0.585 1.975 0.635 2.585 ;
        RECT  0.335 1.275 0.585 1.435 ;
        RECT  0.335 1.975 0.585 2.135 ;
        RECT  0.175 1.275 0.335 2.135 ;
        RECT  0.125 1.515 0.175 2.135 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.510 -0.250 14.720 0.250 ;
        RECT  14.250 -0.250 14.510 1.095 ;
        RECT  13.450 -0.250 14.250 0.250 ;
        RECT  13.190 -0.250 13.450 0.405 ;
        RECT  12.790 -0.250 13.190 0.250 ;
        RECT  12.530 -0.250 12.790 0.405 ;
        RECT  11.670 -0.250 12.530 0.250 ;
        RECT  11.410 -0.250 11.670 0.405 ;
        RECT  10.480 -0.250 11.410 0.250 ;
        RECT  10.220 -0.250 10.480 0.405 ;
        RECT  9.395 -0.250 10.220 0.250 ;
        RECT  9.135 -0.250 9.395 0.405 ;
        RECT  6.645 -0.250 9.135 0.250 ;
        RECT  6.385 -0.250 6.645 0.405 ;
        RECT  4.945 -0.250 6.385 0.250 ;
        RECT  4.685 -0.250 4.945 0.405 ;
        RECT  3.295 -0.250 4.685 0.250 ;
        RECT  3.035 -0.250 3.295 0.405 ;
        RECT  2.205 -0.250 3.035 0.250 ;
        RECT  1.185 -0.250 2.205 0.405 ;
        RECT  0.385 -0.250 1.185 0.250 ;
        RECT  0.125 -0.250 0.385 1.095 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.525 3.440 14.720 3.940 ;
        RECT  14.265 2.255 14.525 3.940 ;
        RECT  13.450 3.440 14.265 3.940 ;
        RECT  13.190 3.285 13.450 3.940 ;
        RECT  11.820 3.440 13.190 3.940 ;
        RECT  11.560 3.285 11.820 3.940 ;
        RECT  10.625 3.440 11.560 3.940 ;
        RECT  10.365 3.285 10.625 3.940 ;
        RECT  9.535 3.440 10.365 3.940 ;
        RECT  9.275 3.285 9.535 3.940 ;
        RECT  6.105 3.440 9.275 3.940 ;
        RECT  5.845 3.285 6.105 3.940 ;
        RECT  4.220 3.440 5.845 3.940 ;
        RECT  3.960 3.065 4.220 3.940 ;
        RECT  2.955 3.440 3.960 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  1.445 3.440 2.695 3.940 ;
        RECT  1.185 3.285 1.445 3.940 ;
        RECT  0.385 3.440 1.185 3.940 ;
        RECT  0.125 2.595 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.560 1.635 13.700 1.795 ;
        RECT  13.400 1.135 13.560 2.115 ;
        RECT  13.050 1.135 13.400 1.295 ;
        RECT  13.050 1.955 13.400 2.115 ;
        RECT  12.610 1.480 13.220 1.740 ;
        RECT  12.790 1.035 13.050 1.295 ;
        RECT  12.790 1.955 13.050 2.555 ;
        RECT  12.450 0.925 12.610 2.770 ;
        RECT  11.430 0.925 12.450 1.085 ;
        RECT  12.270 2.510 12.450 2.770 ;
        RECT  12.110 1.265 12.270 2.325 ;
        RECT  10.970 2.510 12.270 2.670 ;
        RECT  10.890 0.585 12.220 0.745 ;
        RECT  12.010 1.265 12.110 1.645 ;
        RECT  10.790 2.165 12.110 2.325 ;
        RECT  10.450 1.485 12.010 1.645 ;
        RECT  10.450 1.825 11.860 1.985 ;
        RECT  11.170 0.925 11.430 1.305 ;
        RECT  10.730 0.585 10.890 1.175 ;
        RECT  10.630 2.165 10.790 2.765 ;
        RECT  10.630 0.915 10.730 1.175 ;
        RECT  8.755 2.605 10.630 2.765 ;
        RECT  10.290 0.585 10.450 1.645 ;
        RECT  10.290 1.825 10.450 2.425 ;
        RECT  6.155 0.585 10.290 0.745 ;
        RECT  8.595 2.265 10.290 2.425 ;
        RECT  9.055 1.360 9.770 1.520 ;
        RECT  8.895 1.360 9.055 2.055 ;
        RECT  8.855 1.360 8.895 1.520 ;
        RECT  8.795 1.895 8.895 2.055 ;
        RECT  8.695 0.925 8.855 1.520 ;
        RECT  8.595 2.605 8.755 2.880 ;
        RECT  8.595 0.925 8.695 1.185 ;
        RECT  6.985 2.720 8.595 2.880 ;
        RECT  8.255 0.925 8.415 2.540 ;
        RECT  7.295 0.925 8.255 1.085 ;
        RECT  7.325 2.380 8.255 2.540 ;
        RECT  7.915 1.265 8.075 2.200 ;
        RECT  7.045 1.265 7.915 1.425 ;
        RECT  6.935 2.040 7.915 2.200 ;
        RECT  6.495 1.615 7.695 1.775 ;
        RECT  6.885 0.925 7.045 1.425 ;
        RECT  6.825 2.470 6.985 2.880 ;
        RECT  6.675 1.955 6.935 2.215 ;
        RECT  6.785 0.925 6.885 1.175 ;
        RECT  6.335 1.615 6.495 2.425 ;
        RECT  5.015 2.265 6.335 2.425 ;
        RECT  5.995 0.585 6.155 2.085 ;
        RECT  5.835 0.755 5.995 1.015 ;
        RECT  5.265 1.925 5.995 2.085 ;
        RECT  5.265 0.930 5.525 1.190 ;
        RECT  4.915 1.030 5.265 1.190 ;
        RECT  4.915 2.155 5.015 2.425 ;
        RECT  4.755 1.030 4.915 2.425 ;
        RECT  4.305 0.930 4.465 1.935 ;
        RECT  3.650 1.775 4.305 1.935 ;
        RECT  3.625 0.585 3.785 1.255 ;
        RECT  3.390 1.775 3.650 2.375 ;
        RECT  3.390 2.945 3.650 3.205 ;
        RECT  2.495 0.585 3.625 0.745 ;
        RECT  3.275 1.775 3.390 1.935 ;
        RECT  2.245 2.945 3.390 3.105 ;
        RECT  2.185 1.095 3.295 1.255 ;
        RECT  2.085 2.185 2.245 3.105 ;
        RECT  2.025 1.095 2.185 1.345 ;
        RECT  1.675 2.185 2.085 2.345 ;
        RECT  1.675 1.185 2.025 1.345 ;
        RECT  1.235 0.845 1.845 1.005 ;
        RECT  1.585 2.645 1.845 2.905 ;
        RECT  1.515 1.185 1.675 2.345 ;
        RECT  1.235 2.645 1.585 2.805 ;
        RECT  1.415 1.570 1.515 1.830 ;
        RECT  1.075 0.845 1.235 2.805 ;
        RECT  0.805 1.635 1.075 1.795 ;
    END
END BENCX1

MACRO ADDFHX4
    CLASS CORE ;
    FOREIGN ADDFHX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 23.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.265 1.105 23.335 2.045 ;
        RECT  23.040 0.600 23.265 2.045 ;
        RECT  23.030 0.600 23.040 2.920 ;
        RECT  23.005 0.600 23.030 1.200 ;
        RECT  22.780 1.845 23.030 2.920 ;
        END
        ANTENNADIFFAREA     0.8248 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.015 0.540 22.245 1.485 ;
        RECT  21.985 0.540 22.015 2.165 ;
        RECT  21.745 1.290 21.985 2.165 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.575 1.435 20.695 1.725 ;
        RECT  20.365 1.290 20.575 1.725 ;
        RECT  20.340 1.355 20.365 1.725 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.995 1.635 11.410 1.990 ;
        END
        ANTENNAGATEAREA     2.1580 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.500 0.840 1.990 ;
        END
        ANTENNAGATEAREA     0.8086 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  23.775 -0.250 23.920 0.250 ;
        RECT  23.515 -0.250 23.775 1.170 ;
        RECT  22.755 -0.250 23.515 0.250 ;
        RECT  22.495 -0.250 22.755 1.170 ;
        RECT  21.735 -0.250 22.495 0.250 ;
        RECT  21.475 -0.250 21.735 0.755 ;
        RECT  20.795 -0.250 21.475 0.250 ;
        RECT  20.535 -0.250 20.795 0.405 ;
        RECT  19.205 -0.250 20.535 0.250 ;
        RECT  18.945 -0.250 19.205 0.405 ;
        RECT  12.810 -0.250 18.945 0.250 ;
        RECT  12.550 -0.250 12.810 0.405 ;
        RECT  11.670 -0.250 12.550 0.250 ;
        RECT  11.410 -0.250 11.670 0.405 ;
        RECT  3.465 -0.250 11.410 0.250 ;
        RECT  3.205 -0.250 3.465 0.405 ;
        RECT  2.375 -0.250 3.205 0.250 ;
        RECT  2.115 -0.250 2.375 0.405 ;
        RECT  1.435 -0.250 2.115 0.250 ;
        RECT  1.175 -0.250 1.435 0.405 ;
        RECT  0.385 -0.250 1.175 0.250 ;
        RECT  0.125 -0.250 0.385 1.165 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  23.560 3.440 23.920 3.940 ;
        RECT  23.300 2.255 23.560 3.940 ;
        RECT  22.525 3.440 23.300 3.940 ;
        RECT  22.265 2.935 22.525 3.940 ;
        RECT  21.585 3.440 22.265 3.940 ;
        RECT  21.425 2.730 21.585 3.940 ;
        RECT  21.120 2.730 21.425 2.890 ;
        RECT  20.440 3.440 21.425 3.940 ;
        RECT  20.180 3.285 20.440 3.940 ;
        RECT  18.850 3.440 20.180 3.940 ;
        RECT  18.590 3.285 18.850 3.940 ;
        RECT  12.330 3.440 18.590 3.940 ;
        RECT  12.070 2.870 12.330 3.940 ;
        RECT  11.310 3.440 12.070 3.940 ;
        RECT  11.050 2.870 11.310 3.940 ;
        RECT  3.395 3.440 11.050 3.940 ;
        RECT  3.135 2.310 3.395 3.940 ;
        RECT  2.375 3.440 3.135 3.940 ;
        RECT  2.115 2.655 2.375 3.940 ;
        RECT  1.405 3.440 2.115 3.940 ;
        RECT  1.145 3.005 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  22.685 1.405 22.845 1.665 ;
        RECT  22.590 1.505 22.685 1.665 ;
        RECT  22.430 1.505 22.590 2.505 ;
        RECT  20.475 2.345 22.430 2.505 ;
        RECT  21.075 0.950 21.335 1.295 ;
        RECT  20.830 3.100 21.240 3.260 ;
        RECT  20.255 0.950 21.075 1.110 ;
        RECT  20.720 1.905 20.980 2.165 ;
        RECT  20.670 2.945 20.830 3.260 ;
        RECT  20.115 1.905 20.720 2.065 ;
        RECT  15.050 2.945 20.670 3.105 ;
        RECT  20.315 2.345 20.475 2.765 ;
        RECT  17.800 2.605 20.315 2.765 ;
        RECT  20.115 0.495 20.255 1.110 ;
        RECT  19.995 0.495 20.115 2.065 ;
        RECT  19.955 0.590 19.995 2.065 ;
        RECT  17.245 0.590 19.955 0.750 ;
        RECT  19.900 1.825 19.955 2.065 ;
        RECT  19.640 1.825 19.900 2.215 ;
        RECT  19.485 0.930 19.745 1.190 ;
        RECT  18.790 1.825 19.640 1.985 ;
        RECT  18.665 0.930 19.485 1.090 ;
        RECT  18.325 2.265 19.390 2.425 ;
        RECT  18.565 0.930 18.665 1.190 ;
        RECT  18.405 0.930 18.565 1.545 ;
        RECT  17.615 1.385 18.405 1.545 ;
        RECT  18.050 2.165 18.325 2.425 ;
        RECT  17.895 0.945 18.155 1.205 ;
        RECT  17.210 2.165 18.050 2.325 ;
        RECT  16.870 0.945 17.895 1.105 ;
        RECT  17.540 2.505 17.800 2.765 ;
        RECT  17.355 1.285 17.615 1.545 ;
        RECT  16.870 2.605 17.540 2.765 ;
        RECT  17.210 1.385 17.355 1.545 ;
        RECT  16.985 0.590 17.245 0.765 ;
        RECT  17.050 1.385 17.210 2.425 ;
        RECT  16.195 0.590 16.985 0.750 ;
        RECT  16.710 0.945 16.870 2.765 ;
        RECT  16.445 0.945 16.710 1.205 ;
        RECT  15.810 2.605 16.710 2.765 ;
        RECT  16.370 2.105 16.530 2.425 ;
        RECT  15.560 2.265 16.370 2.425 ;
        RECT  16.095 0.590 16.195 1.135 ;
        RECT  15.935 0.555 16.095 1.715 ;
        RECT  15.245 0.555 15.935 0.715 ;
        RECT  15.560 1.555 15.935 1.715 ;
        RECT  15.585 0.895 15.685 1.155 ;
        RECT  15.425 0.895 15.585 1.375 ;
        RECT  15.400 1.555 15.560 2.425 ;
        RECT  14.150 1.215 15.425 1.375 ;
        RECT  15.300 2.105 15.400 2.425 ;
        RECT  14.490 2.265 15.300 2.425 ;
        RECT  15.085 0.555 15.245 0.980 ;
        RECT  14.905 0.820 15.085 0.980 ;
        RECT  14.790 2.695 15.050 3.105 ;
        RECT  14.645 0.430 14.905 0.640 ;
        RECT  14.150 2.945 14.790 3.105 ;
        RECT  13.310 0.480 14.645 0.640 ;
        RECT  13.660 0.820 14.645 0.980 ;
        RECT  14.330 2.060 14.490 2.660 ;
        RECT  14.100 1.215 14.150 3.105 ;
        RECT  13.990 1.160 14.100 3.105 ;
        RECT  13.840 1.160 13.990 1.375 ;
        RECT  13.350 2.945 13.990 3.105 ;
        RECT  13.660 1.555 13.810 2.635 ;
        RECT  13.650 0.820 13.660 2.635 ;
        RECT  13.500 0.820 13.650 1.715 ;
        RECT  12.825 2.355 13.650 2.515 ;
        RECT  13.100 0.925 13.500 1.085 ;
        RECT  13.320 1.900 13.440 2.160 ;
        RECT  13.090 2.845 13.350 3.105 ;
        RECT  13.160 1.265 13.320 2.160 ;
        RECT  13.150 0.480 13.310 0.745 ;
        RECT  12.920 1.265 13.160 1.425 ;
        RECT  12.920 0.585 13.150 0.745 ;
        RECT  12.580 1.635 12.980 1.795 ;
        RECT  12.760 0.585 12.920 1.425 ;
        RECT  12.580 2.355 12.825 3.065 ;
        RECT  8.655 0.585 12.760 0.745 ;
        RECT  12.420 0.925 12.580 1.795 ;
        RECT  11.950 2.355 12.580 2.515 ;
        RECT  8.995 0.925 12.420 1.085 ;
        RECT  11.950 1.265 12.240 1.425 ;
        RECT  11.820 1.265 11.950 2.515 ;
        RECT  11.790 1.265 11.820 3.130 ;
        RECT  10.835 1.265 11.790 1.425 ;
        RECT  11.560 2.350 11.790 3.130 ;
        RECT  10.710 2.350 11.560 2.515 ;
        RECT  10.610 2.350 10.710 3.195 ;
        RECT  10.450 1.900 10.610 3.195 ;
        RECT  10.270 1.265 10.525 1.425 ;
        RECT  10.110 1.265 10.270 3.220 ;
        RECT  9.335 1.265 10.110 1.425 ;
        RECT  4.925 3.060 10.110 3.220 ;
        RECT  9.770 1.725 9.930 2.880 ;
        RECT  8.995 1.725 9.770 1.885 ;
        RECT  6.455 2.720 9.770 2.880 ;
        RECT  9.430 2.250 9.590 2.540 ;
        RECT  8.560 2.380 9.430 2.540 ;
        RECT  9.175 1.265 9.335 1.525 ;
        RECT  8.835 0.925 8.995 1.885 ;
        RECT  8.560 0.585 8.655 1.075 ;
        RECT  8.400 0.585 8.560 2.540 ;
        RECT  8.395 0.585 8.400 1.075 ;
        RECT  8.300 2.280 8.400 2.540 ;
        RECT  7.635 0.585 8.395 0.745 ;
        RECT  7.475 2.380 8.300 2.540 ;
        RECT  8.045 0.955 8.145 1.215 ;
        RECT  7.885 0.955 8.045 2.200 ;
        RECT  7.760 1.730 7.885 2.200 ;
        RECT  7.030 1.730 7.760 1.890 ;
        RECT  7.375 0.585 7.635 1.205 ;
        RECT  7.215 2.280 7.475 2.540 ;
        RECT  7.030 0.855 7.125 1.115 ;
        RECT  7.025 0.855 7.030 1.890 ;
        RECT  6.865 0.585 7.025 1.890 ;
        RECT  6.865 2.175 6.965 2.435 ;
        RECT  6.105 0.585 6.865 0.745 ;
        RECT  6.705 1.730 6.865 2.435 ;
        RECT  5.945 1.730 6.705 1.890 ;
        RECT  6.565 0.930 6.615 1.190 ;
        RECT  6.355 0.930 6.565 1.290 ;
        RECT  6.195 2.175 6.455 2.880 ;
        RECT  5.595 1.125 6.355 1.290 ;
        RECT  5.435 2.720 6.195 2.880 ;
        RECT  5.845 0.585 6.105 0.945 ;
        RECT  5.785 1.730 5.945 2.435 ;
        RECT  0.895 0.585 5.845 0.745 ;
        RECT  5.685 2.175 5.785 2.435 ;
        RECT  5.495 0.965 5.595 1.290 ;
        RECT  5.335 0.965 5.495 1.425 ;
        RECT  5.385 2.280 5.435 2.880 ;
        RECT  5.175 2.105 5.385 2.880 ;
        RECT  4.445 1.265 5.335 1.425 ;
        RECT  4.445 2.105 5.175 2.265 ;
        RECT  4.005 0.925 5.085 1.085 ;
        RECT  4.665 2.445 4.925 3.220 ;
        RECT  3.905 3.060 4.665 3.220 ;
        RECT  4.415 1.265 4.445 2.265 ;
        RECT  4.285 1.265 4.415 2.740 ;
        RECT  4.155 2.105 4.285 2.740 ;
        RECT  3.905 0.925 4.005 1.185 ;
        RECT  3.745 0.925 3.905 3.220 ;
        RECT  2.925 1.025 3.745 1.185 ;
        RECT  3.650 1.965 3.745 3.220 ;
        RECT  3.645 1.965 3.650 3.080 ;
        RECT  2.885 1.965 3.645 2.125 ;
        RECT  2.665 0.925 2.925 1.185 ;
        RECT  2.625 1.965 2.885 2.905 ;
        RECT  1.975 1.580 2.160 1.840 ;
        RECT  1.815 1.035 1.975 2.215 ;
        RECT  1.715 1.035 1.815 1.295 ;
        RECT  1.715 1.955 1.815 2.215 ;
        RECT  1.025 1.025 1.185 2.330 ;
        RECT  0.895 1.025 1.025 1.185 ;
        RECT  0.895 2.170 1.025 2.330 ;
        RECT  0.635 0.585 0.895 1.185 ;
        RECT  0.635 2.170 0.895 3.110 ;
    END
END ADDFHX4

MACRO ADDFHX2
    CLASS CORE ;
    FOREIGN ADDFHX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.385 0.695 14.595 2.920 ;
        RECT  14.335 0.695 14.385 1.295 ;
        RECT  14.335 1.980 14.385 2.920 ;
        END
        ANTENNADIFFAREA     0.7528 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.575 1.515 13.675 1.990 ;
        RECT  13.415 0.495 13.575 2.225 ;
        RECT  13.315 0.495 13.415 0.755 ;
        RECT  13.335 1.965 13.415 2.225 ;
        END
        ANTENNADIFFAREA     0.5551 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 1.500 12.795 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.235 1.635 8.650 1.990 ;
        RECT  8.195 1.635 8.235 1.795 ;
        END
        ANTENNAGATEAREA     1.0868 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.500 0.380 1.990 ;
        END
        ANTENNAGATEAREA     0.4030 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.085 -0.250 14.720 0.250 ;
        RECT  13.825 -0.250 14.085 1.170 ;
        RECT  12.595 -0.250 13.825 0.250 ;
        RECT  12.335 -0.250 12.595 0.405 ;
        RECT  9.235 -0.250 12.335 0.250 ;
        RECT  8.975 -0.250 9.235 0.405 ;
        RECT  2.235 -0.250 8.975 0.250 ;
        RECT  1.975 -0.250 2.235 0.405 ;
        RECT  0.925 -0.250 1.975 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.060 3.440 14.720 3.940 ;
        RECT  13.800 2.945 14.060 3.940 ;
        RECT  12.490 3.440 13.800 3.940 ;
        RECT  12.230 3.285 12.490 3.940 ;
        RECT  8.825 3.440 12.230 3.940 ;
        RECT  8.565 2.870 8.825 3.940 ;
        RECT  2.125 3.440 8.565 3.940 ;
        RECT  1.865 2.935 2.125 3.940 ;
        RECT  0.895 3.440 1.865 3.940 ;
        RECT  0.635 2.955 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.125 1.570 14.175 1.830 ;
        RECT  14.015 1.570 14.125 2.760 ;
        RECT  13.965 1.575 14.015 2.760 ;
        RECT  11.455 2.600 13.965 2.760 ;
        RECT  10.540 2.945 13.290 3.105 ;
        RECT  12.910 1.035 13.170 1.295 ;
        RECT  12.310 2.170 13.035 2.330 ;
        RECT  12.310 1.135 12.910 1.295 ;
        RECT  12.150 0.695 12.310 2.330 ;
        RECT  11.000 0.695 12.150 0.855 ;
        RECT  11.975 1.810 12.150 2.080 ;
        RECT  11.810 1.035 11.970 1.630 ;
        RECT  11.795 2.260 11.950 2.420 ;
        RECT  11.795 1.470 11.810 1.630 ;
        RECT  11.635 1.470 11.795 2.420 ;
        RECT  11.455 1.035 11.510 1.295 ;
        RECT  11.295 1.035 11.455 2.760 ;
        RECT  11.250 1.035 11.295 1.295 ;
        RECT  11.180 2.500 11.295 2.760 ;
        RECT  10.880 0.695 11.000 1.220 ;
        RECT  10.840 0.695 10.880 2.665 ;
        RECT  10.720 0.960 10.840 2.665 ;
        RECT  10.400 0.430 10.660 0.745 ;
        RECT  10.380 0.925 10.540 3.105 ;
        RECT  9.350 0.585 10.400 0.745 ;
        RECT  10.230 0.925 10.380 1.085 ;
        RECT  9.735 2.695 10.380 2.955 ;
        RECT  10.040 1.545 10.200 2.515 ;
        RECT  10.025 1.545 10.040 1.705 ;
        RECT  9.320 2.355 10.040 2.515 ;
        RECT  9.865 0.925 10.025 1.705 ;
        RECT  9.530 0.925 9.865 1.085 ;
        RECT  9.700 1.905 9.860 2.165 ;
        RECT  9.685 1.905 9.700 2.065 ;
        RECT  9.525 1.265 9.685 2.065 ;
        RECT  9.350 1.265 9.525 1.425 ;
        RECT  9.190 0.585 9.350 1.425 ;
        RECT  9.010 1.635 9.345 1.795 ;
        RECT  9.075 2.355 9.320 3.065 ;
        RECT  6.675 0.585 9.190 0.745 ;
        RECT  8.315 2.355 9.075 2.515 ;
        RECT  8.850 0.925 9.010 1.795 ;
        RECT  7.015 0.925 8.850 1.085 ;
        RECT  8.005 1.265 8.665 1.425 ;
        RECT  8.055 2.355 8.315 3.130 ;
        RECT  8.005 2.355 8.055 2.515 ;
        RECT  7.845 1.265 8.005 2.515 ;
        RECT  7.505 1.270 7.665 3.190 ;
        RECT  7.220 1.270 7.505 1.430 ;
        RECT  3.655 3.030 7.505 3.190 ;
        RECT  7.165 1.675 7.325 2.850 ;
        RECT  7.015 1.675 7.165 1.835 ;
        RECT  4.565 2.690 7.165 2.850 ;
        RECT  6.855 0.925 7.015 1.835 ;
        RECT  6.675 2.250 6.985 2.510 ;
        RECT  6.515 0.585 6.675 2.510 ;
        RECT  5.825 0.585 6.515 0.745 ;
        RECT  5.585 2.350 6.515 2.510 ;
        RECT  6.230 0.960 6.335 1.220 ;
        RECT  6.125 0.960 6.230 2.055 ;
        RECT  6.075 0.960 6.125 2.165 ;
        RECT  6.070 1.010 6.075 2.165 ;
        RECT  5.850 1.895 6.070 2.165 ;
        RECT  5.210 1.895 5.850 2.055 ;
        RECT  5.650 0.585 5.825 1.150 ;
        RECT  5.565 0.890 5.650 1.150 ;
        RECT  5.325 2.250 5.585 2.510 ;
        RECT  5.210 0.920 5.315 1.180 ;
        RECT  5.205 0.920 5.210 2.055 ;
        RECT  5.075 0.585 5.205 2.055 ;
        RECT  5.045 0.585 5.075 2.435 ;
        RECT  4.265 0.585 5.045 0.745 ;
        RECT  4.815 1.895 5.045 2.435 ;
        RECT  4.055 1.895 4.815 2.055 ;
        RECT  4.705 0.930 4.805 1.190 ;
        RECT  4.545 0.930 4.705 1.530 ;
        RECT  4.305 2.250 4.565 2.850 ;
        RECT  3.325 1.370 4.545 1.530 ;
        RECT  3.165 2.590 4.305 2.750 ;
        RECT  4.005 0.470 4.265 0.745 ;
        RECT  3.895 1.895 4.055 2.380 ;
        RECT  0.725 0.585 4.005 0.745 ;
        RECT  3.795 2.220 3.895 2.380 ;
        RECT  3.605 0.960 3.865 1.190 ;
        RECT  3.395 2.930 3.655 3.190 ;
        RECT  2.785 0.960 3.605 1.120 ;
        RECT  2.635 3.030 3.395 3.190 ;
        RECT  3.165 1.300 3.325 1.530 ;
        RECT  3.065 1.300 3.165 2.750 ;
        RECT  3.005 1.365 3.065 2.750 ;
        RECT  2.885 2.490 3.005 2.750 ;
        RECT  2.525 0.960 2.785 1.235 ;
        RECT  2.375 2.575 2.635 3.190 ;
        RECT  1.835 1.075 2.525 1.235 ;
        RECT  1.805 2.575 2.375 2.735 ;
        RECT  1.805 0.975 1.835 1.235 ;
        RECT  1.645 0.975 1.805 2.735 ;
        RECT  1.575 0.975 1.645 1.235 ;
        RECT  1.615 2.575 1.645 2.735 ;
        RECT  1.455 2.575 1.615 3.005 ;
        RECT  1.325 1.585 1.465 1.845 ;
        RECT  1.355 2.745 1.455 3.005 ;
        RECT  1.155 1.035 1.325 2.215 ;
        RECT  1.065 1.035 1.155 1.295 ;
        RECT  1.065 1.955 1.155 2.215 ;
        RECT  0.565 0.585 0.725 2.330 ;
        RECT  0.385 0.585 0.565 0.745 ;
        RECT  0.385 2.170 0.565 2.330 ;
        RECT  0.125 0.585 0.385 1.185 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END ADDFHX2

MACRO ADDFHX1
    CLASS CORE ;
    FOREIGN ADDFHX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.245 0.985 10.455 2.215 ;
        RECT  10.195 0.985 10.245 1.355 ;
        RECT  10.195 1.925 10.245 2.215 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.505 1.105 9.535 1.990 ;
        RECT  9.395 0.955 9.505 1.990 ;
        RECT  9.210 0.955 9.395 2.215 ;
        RECT  9.135 1.955 9.210 2.215 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.360 1.555 8.615 2.080 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.725 1.290 4.935 1.915 ;
        RECT  4.695 1.655 4.725 1.915 ;
        END
        ANTENNAGATEAREA     0.5382 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.500 0.380 1.990 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.055 -0.250 10.580 0.250 ;
        RECT  9.795 -0.250 10.055 0.405 ;
        RECT  8.445 -0.250 9.795 0.250 ;
        RECT  8.185 -0.250 8.445 0.405 ;
        RECT  5.275 -0.250 8.185 0.250 ;
        RECT  5.015 -0.250 5.275 0.405 ;
        RECT  1.620 -0.250 5.015 0.250 ;
        RECT  0.680 -0.250 1.620 0.405 ;
        RECT  0.000 -0.250 0.680 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.945 3.440 10.580 3.940 ;
        RECT  9.685 3.285 9.945 3.940 ;
        RECT  8.175 3.440 9.685 3.940 ;
        RECT  7.915 3.285 8.175 3.940 ;
        RECT  4.745 3.440 7.915 3.940 ;
        RECT  4.485 2.870 4.745 3.940 ;
        RECT  1.280 3.440 4.485 3.940 ;
        RECT  1.020 2.790 1.280 3.940 ;
        RECT  0.000 3.440 1.020 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.025 2.605 10.285 2.925 ;
        RECT  7.315 2.605 10.025 2.765 ;
        RECT  6.365 2.945 9.515 3.105 ;
        RECT  8.955 0.955 8.995 1.215 ;
        RECT  8.895 0.955 8.955 2.425 ;
        RECT  8.795 0.610 8.895 2.425 ;
        RECT  8.735 0.610 8.795 1.215 ;
        RECT  8.140 2.265 8.795 2.425 ;
        RECT  6.975 0.610 8.735 0.770 ;
        RECT  7.995 1.925 8.140 2.425 ;
        RECT  7.945 0.960 8.045 1.220 ;
        RECT  7.980 1.825 7.995 2.425 ;
        RECT  7.835 1.825 7.980 2.085 ;
        RECT  7.785 0.960 7.945 1.640 ;
        RECT  7.655 1.480 7.785 1.640 ;
        RECT  7.655 2.265 7.775 2.425 ;
        RECT  7.495 1.480 7.655 2.425 ;
        RECT  7.315 0.960 7.535 1.220 ;
        RECT  7.275 0.960 7.315 2.765 ;
        RECT  7.155 1.060 7.275 2.765 ;
        RECT  7.005 2.345 7.155 2.605 ;
        RECT  6.815 0.610 6.975 1.255 ;
        RECT  6.810 1.095 6.815 1.255 ;
        RECT  6.705 1.095 6.810 2.595 ;
        RECT  6.650 1.095 6.705 2.665 ;
        RECT  6.545 2.405 6.650 2.665 ;
        RECT  6.445 0.475 6.605 0.745 ;
        RECT  6.365 0.950 6.465 2.115 ;
        RECT  5.615 0.585 6.445 0.745 ;
        RECT  6.305 0.950 6.365 3.105 ;
        RECT  6.205 1.955 6.305 3.105 ;
        RECT  5.720 2.945 6.205 3.105 ;
        RECT  5.865 0.945 6.025 2.755 ;
        RECT  5.795 0.945 5.865 1.205 ;
        RECT  5.240 2.595 5.865 2.755 ;
        RECT  5.615 1.385 5.685 2.415 ;
        RECT  5.525 0.585 5.615 2.415 ;
        RECT  5.455 0.585 5.525 1.545 ;
        RECT  5.425 2.255 5.525 2.415 ;
        RECT  3.835 0.585 5.455 0.745 ;
        RECT  5.275 1.725 5.345 1.985 ;
        RECT  5.115 0.925 5.275 1.985 ;
        RECT  4.995 2.425 5.240 3.025 ;
        RECT  4.175 0.925 5.115 1.085 ;
        RECT  4.435 2.425 4.995 2.585 ;
        RECT  4.355 1.265 4.515 2.125 ;
        RECT  4.275 2.305 4.435 2.585 ;
        RECT  4.095 1.965 4.355 2.125 ;
        RECT  4.015 0.925 4.175 1.785 ;
        RECT  3.935 1.965 4.095 3.190 ;
        RECT  3.755 1.625 4.015 1.785 ;
        RECT  1.995 3.030 3.935 3.190 ;
        RECT  3.675 0.585 3.835 1.445 ;
        RECT  3.595 1.625 3.755 2.850 ;
        RECT  3.415 1.285 3.675 1.445 ;
        RECT  2.435 2.690 3.595 2.850 ;
        RECT  3.255 1.285 3.415 2.510 ;
        RECT  3.075 0.845 3.375 1.105 ;
        RECT  2.945 0.585 3.075 1.885 ;
        RECT  2.915 0.585 2.945 2.510 ;
        RECT  0.725 0.585 2.915 0.745 ;
        RECT  2.785 1.725 2.915 2.510 ;
        RECT  2.685 2.250 2.785 2.510 ;
        RECT  2.575 1.015 2.735 1.530 ;
        RECT  2.435 1.370 2.575 1.530 ;
        RECT  2.275 1.370 2.435 2.850 ;
        RECT  2.015 0.925 2.275 1.185 ;
        RECT  2.175 2.250 2.275 2.850 ;
        RECT  1.995 1.025 2.015 1.185 ;
        RECT  1.835 1.025 1.995 3.190 ;
        RECT  1.665 2.675 1.835 2.935 ;
        RECT  1.365 1.585 1.475 1.845 ;
        RECT  1.335 1.035 1.365 1.845 ;
        RECT  1.175 1.035 1.335 2.215 ;
        RECT  1.105 1.035 1.175 1.295 ;
        RECT  1.075 1.955 1.175 2.215 ;
        RECT  0.565 0.585 0.725 2.330 ;
        RECT  0.125 1.035 0.565 1.295 ;
        RECT  0.385 2.170 0.565 2.330 ;
        RECT  0.125 2.170 0.385 2.430 ;
    END
END ADDFHX1

MACRO ADDFHXL
    CLASS CORE ;
    FOREIGN ADDFHXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.985 1.105 9.995 2.375 ;
        RECT  9.785 1.035 9.985 2.375 ;
        RECT  9.725 1.035 9.785 1.355 ;
        RECT  9.735 2.115 9.785 2.375 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.070 1.925 9.075 2.400 ;
        RECT  8.910 0.610 9.070 2.400 ;
        RECT  8.835 0.610 8.910 0.770 ;
        RECT  8.865 1.925 8.910 2.400 ;
        RECT  8.835 2.115 8.865 2.375 ;
        RECT  8.575 0.510 8.835 0.770 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.155 1.735 8.275 1.995 ;
        RECT  7.995 1.290 8.155 1.995 ;
        RECT  7.945 1.290 7.995 1.580 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.170 1.290 4.475 1.795 ;
        END
        ANTENNAGATEAREA     0.2496 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.480 0.795 1.990 ;
        RECT  0.495 1.480 0.585 1.740 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.405 -0.250 10.120 0.250 ;
        RECT  9.145 -0.250 9.405 0.405 ;
        RECT  8.145 -0.250 9.145 0.250 ;
        RECT  7.885 -0.250 8.145 0.405 ;
        RECT  5.095 -0.250 7.885 0.250 ;
        RECT  4.835 -0.250 5.095 0.405 ;
        RECT  1.220 -0.250 4.835 0.250 ;
        RECT  0.960 -0.250 1.220 0.405 ;
        RECT  0.000 -0.250 0.960 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.595 3.440 10.120 3.940 ;
        RECT  9.335 3.285 9.595 3.940 ;
        RECT  7.985 3.440 9.335 3.940 ;
        RECT  7.725 3.285 7.985 3.940 ;
        RECT  4.285 3.440 7.725 3.940 ;
        RECT  4.025 2.815 4.285 3.940 ;
        RECT  0.490 3.440 4.025 3.940 ;
        RECT  0.230 3.285 0.490 3.940 ;
        RECT  0.000 3.440 0.230 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.865 2.605 9.825 2.765 ;
        RECT  5.965 2.945 9.215 3.105 ;
        RECT  8.625 1.030 8.725 1.290 ;
        RECT  8.615 0.950 8.625 1.290 ;
        RECT  8.455 0.950 8.615 2.425 ;
        RECT  8.235 0.950 8.455 1.110 ;
        RECT  7.795 2.265 8.455 2.425 ;
        RECT  8.075 0.610 8.235 1.110 ;
        RECT  6.645 0.610 8.075 0.770 ;
        RECT  7.635 1.825 7.795 2.425 ;
        RECT  7.615 1.030 7.715 1.290 ;
        RECT  7.455 1.030 7.615 1.645 ;
        RECT  7.295 1.485 7.455 2.425 ;
        RECT  7.145 2.265 7.295 2.425 ;
        RECT  7.115 1.025 7.155 1.290 ;
        RECT  6.955 1.025 7.115 2.070 ;
        RECT  6.865 1.910 6.955 2.070 ;
        RECT  6.705 1.910 6.865 2.765 ;
        RECT  6.605 2.605 6.705 2.765 ;
        RECT  6.485 0.610 6.645 1.720 ;
        RECT  6.305 1.560 6.485 1.720 ;
        RECT  6.145 0.510 6.305 0.770 ;
        RECT  6.145 1.560 6.305 2.765 ;
        RECT  5.965 1.080 6.185 1.240 ;
        RECT  5.285 0.585 6.145 0.745 ;
        RECT  5.805 1.080 5.965 3.105 ;
        RECT  5.165 2.930 5.805 3.105 ;
        RECT  5.465 1.030 5.625 2.750 ;
        RECT  4.885 2.590 5.465 2.750 ;
        RECT  5.125 0.585 5.285 2.410 ;
        RECT  3.130 0.585 5.125 0.745 ;
        RECT  4.805 2.250 5.125 2.410 ;
        RECT  4.815 1.720 4.945 1.985 ;
        RECT  4.625 2.590 4.885 2.870 ;
        RECT  4.655 0.925 4.815 1.985 ;
        RECT  3.470 0.925 4.655 1.085 ;
        RECT  4.465 2.405 4.625 2.750 ;
        RECT  4.155 2.405 4.465 2.565 ;
        RECT  3.995 2.140 4.155 2.565 ;
        RECT  3.650 1.265 3.810 2.385 ;
        RECT  3.620 2.225 3.650 2.385 ;
        RECT  3.460 2.225 3.620 3.190 ;
        RECT  3.310 0.925 3.470 2.045 ;
        RECT  1.480 3.030 3.460 3.190 ;
        RECT  3.280 1.885 3.310 2.045 ;
        RECT  3.120 1.885 3.280 2.850 ;
        RECT  2.970 0.585 3.130 1.700 ;
        RECT  1.920 2.690 3.120 2.850 ;
        RECT  2.815 1.540 2.970 1.700 ;
        RECT  2.815 2.350 2.940 2.510 ;
        RECT  2.655 1.540 2.815 2.510 ;
        RECT  2.475 1.035 2.670 1.295 ;
        RECT  2.315 0.695 2.475 2.510 ;
        RECT  0.640 0.695 2.315 0.855 ;
        RECT  2.170 2.350 2.315 2.510 ;
        RECT  1.950 1.035 2.110 1.795 ;
        RECT  1.920 1.635 1.950 1.795 ;
        RECT  1.760 1.635 1.920 2.850 ;
        RECT  1.660 2.390 1.760 2.650 ;
        RECT  1.480 1.035 1.650 1.295 ;
        RECT  1.320 1.035 1.480 3.190 ;
        RECT  1.150 2.510 1.320 2.670 ;
        RECT  0.975 1.135 1.135 2.330 ;
        RECT  0.590 1.135 0.975 1.295 ;
        RECT  0.855 2.170 0.975 2.330 ;
        RECT  0.695 2.170 0.855 2.625 ;
        RECT  0.385 2.465 0.695 2.625 ;
        RECT  0.380 0.525 0.640 0.855 ;
        RECT  0.430 1.035 0.590 1.295 ;
        RECT  0.285 1.955 0.385 2.215 ;
        RECT  0.125 2.465 0.385 2.725 ;
        RECT  0.250 0.695 0.380 0.855 ;
        RECT  0.250 1.475 0.285 2.215 ;
        RECT  0.125 0.695 0.250 2.215 ;
        RECT  0.090 0.695 0.125 1.635 ;
    END
END ADDFHXL

MACRO ADDFX4
    CLASS CORE ;
    FOREIGN ADDFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.945 1.095 9.995 2.585 ;
        RECT  9.765 0.695 9.945 2.945 ;
        RECT  9.685 0.695 9.765 1.295 ;
        RECT  9.685 2.005 9.765 2.945 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.665 0.695 8.925 1.295 ;
        RECT  8.615 1.960 8.925 2.220 ;
        RECT  8.615 0.880 8.665 1.295 ;
        RECT  8.590 0.880 8.615 2.220 ;
        RECT  8.355 1.035 8.590 2.220 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 2.260 6.320 2.520 ;
        RECT  6.265 1.700 6.315 2.520 ;
        RECT  6.105 1.310 6.265 2.520 ;
        RECT  6.100 1.310 6.105 1.925 ;
        RECT  6.060 2.260 6.105 2.520 ;
        END
        ANTENNAGATEAREA     0.1976 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.490 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.510 3.165 1.990 ;
        RECT  2.645 1.510 2.885 1.825 ;
        END
        ANTENNAGATEAREA     0.2769 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.455 -0.250 10.580 0.250 ;
        RECT  10.195 -0.250 10.455 1.095 ;
        RECT  9.435 -0.250 10.195 0.250 ;
        RECT  9.175 -0.250 9.435 1.095 ;
        RECT  8.385 -0.250 9.175 0.250 ;
        RECT  8.125 -0.250 8.385 0.405 ;
        RECT  6.570 -0.250 8.125 0.250 ;
        RECT  6.310 -0.250 6.570 0.405 ;
        RECT  3.115 -0.250 6.310 0.250 ;
        RECT  2.855 -0.250 3.115 0.575 ;
        RECT  0.925 -0.250 2.855 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.455 3.440 10.580 3.940 ;
        RECT  10.195 2.255 10.455 3.940 ;
        RECT  9.435 3.440 10.195 3.940 ;
        RECT  9.175 2.935 9.435 3.940 ;
        RECT  8.420 3.440 9.175 3.940 ;
        RECT  8.160 2.895 8.420 3.940 ;
        RECT  8.125 3.285 8.160 3.940 ;
        RECT  6.420 3.440 8.125 3.940 ;
        RECT  6.160 3.285 6.420 3.940 ;
        RECT  3.155 3.440 6.160 3.940 ;
        RECT  2.895 3.285 3.155 3.940 ;
        RECT  0.925 3.440 2.895 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.475 1.565 9.575 1.825 ;
        RECT  9.315 1.565 9.475 2.690 ;
        RECT  7.330 2.530 9.315 2.690 ;
        RECT  6.760 2.870 7.980 3.030 ;
        RECT  7.820 1.035 7.940 1.295 ;
        RECT  7.820 2.090 7.870 2.350 ;
        RECT  7.660 0.615 7.820 2.350 ;
        RECT  6.130 0.615 7.660 0.775 ;
        RECT  7.610 2.090 7.660 2.350 ;
        RECT  7.330 1.035 7.430 1.295 ;
        RECT  7.170 1.035 7.330 2.690 ;
        RECT  7.120 2.280 7.170 2.690 ;
        RECT  7.070 2.280 7.120 2.540 ;
        RECT  6.720 1.035 6.920 1.295 ;
        RECT  6.720 2.125 6.820 2.385 ;
        RECT  6.600 2.735 6.760 3.030 ;
        RECT  6.560 0.955 6.720 2.385 ;
        RECT  5.450 2.735 6.600 2.895 ;
        RECT  5.790 0.955 6.560 1.115 ;
        RECT  5.970 0.530 6.130 0.775 ;
        RECT  4.050 0.530 5.970 0.690 ;
        RECT  5.790 1.295 5.920 1.455 ;
        RECT  5.630 0.885 5.790 1.115 ;
        RECT  5.630 1.295 5.790 2.545 ;
        RECT  4.480 0.885 5.630 1.045 ;
        RECT  5.290 1.275 5.450 2.895 ;
        RECT  5.120 1.275 5.290 1.435 ;
        RECT  4.810 2.735 5.290 2.895 ;
        RECT  4.950 1.615 5.110 2.555 ;
        RECT  4.820 1.615 4.950 1.775 ;
        RECT  4.560 2.395 4.950 2.555 ;
        RECT  4.660 1.225 4.820 1.775 ;
        RECT  4.480 1.955 4.770 2.215 ;
        RECT  4.460 2.395 4.560 2.795 ;
        RECT  4.320 0.885 4.480 2.215 ;
        RECT  4.400 2.395 4.460 3.010 ;
        RECT  4.300 2.535 4.400 3.010 ;
        RECT  4.050 2.055 4.320 2.215 ;
        RECT  2.320 2.850 4.300 3.010 ;
        RECT  3.540 1.485 4.140 1.745 ;
        RECT  3.890 0.530 4.050 1.305 ;
        RECT  3.950 2.055 4.050 2.425 ;
        RECT  3.840 2.055 3.950 2.670 ;
        RECT  3.790 0.755 3.890 1.305 ;
        RECT  3.790 2.165 3.840 2.670 ;
        RECT  2.530 0.755 3.790 0.915 ;
        RECT  2.320 2.510 3.790 2.670 ;
        RECT  3.380 1.095 3.540 2.330 ;
        RECT  2.305 1.095 3.380 1.255 ;
        RECT  2.660 2.170 3.380 2.330 ;
        RECT  2.500 2.015 2.660 2.330 ;
        RECT  2.370 0.695 2.530 0.915 ;
        RECT  2.355 2.015 2.500 2.175 ;
        RECT  1.665 0.695 2.370 0.855 ;
        RECT  2.175 2.380 2.320 2.670 ;
        RECT  2.160 2.850 2.320 3.260 ;
        RECT  2.160 1.595 2.175 2.670 ;
        RECT  2.015 1.595 2.160 2.540 ;
        RECT  1.495 3.100 2.160 3.260 ;
        RECT  2.005 1.595 2.015 1.755 ;
        RECT  1.845 1.045 2.005 1.755 ;
        RECT  1.835 2.760 1.980 2.920 ;
        RECT  1.665 1.965 1.835 2.225 ;
        RECT  1.675 2.480 1.835 2.920 ;
        RECT  1.325 2.480 1.675 2.640 ;
        RECT  1.505 0.695 1.665 2.225 ;
        RECT  1.335 2.945 1.495 3.260 ;
        RECT  0.385 2.945 1.335 3.105 ;
        RECT  1.165 1.035 1.325 2.640 ;
        RECT  1.075 1.035 1.165 1.295 ;
        RECT  1.065 2.070 1.165 2.640 ;
        RECT  0.745 1.500 0.985 1.760 ;
        RECT  0.585 1.135 0.745 2.330 ;
        RECT  0.385 1.135 0.585 1.295 ;
        RECT  0.385 2.170 0.585 2.330 ;
        RECT  0.125 0.695 0.385 1.295 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END ADDFX4

MACRO ADDFX2
    CLASS CORE ;
    FOREIGN ADDFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.325 0.695 9.535 2.945 ;
        RECT  9.275 0.695 9.325 1.295 ;
        RECT  9.275 2.005 9.325 2.945 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.455 1.515 8.615 1.990 ;
        RECT  8.450 1.135 8.455 2.265 ;
        RECT  8.295 0.695 8.450 2.265 ;
        RECT  8.190 0.695 8.295 1.295 ;
        RECT  8.195 2.005 8.295 2.265 ;
        END
        ANTENNADIFFAREA     0.7195 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 2.260 6.320 2.520 ;
        RECT  6.265 1.700 6.315 2.520 ;
        RECT  6.105 1.310 6.265 2.520 ;
        RECT  6.100 1.310 6.105 1.925 ;
        RECT  6.060 2.260 6.105 2.520 ;
        END
        ANTENNAGATEAREA     0.1976 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.490 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.510 3.165 1.990 ;
        RECT  2.645 1.510 2.885 1.825 ;
        END
        ANTENNAGATEAREA     0.2769 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.995 -0.250 9.660 0.250 ;
        RECT  8.735 -0.250 8.995 1.145 ;
        RECT  6.570 -0.250 8.735 0.250 ;
        RECT  6.310 -0.250 6.570 0.405 ;
        RECT  3.115 -0.250 6.310 0.250 ;
        RECT  2.855 -0.250 3.115 0.575 ;
        RECT  0.925 -0.250 2.855 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.995 3.440 9.660 3.940 ;
        RECT  8.735 2.880 8.995 3.940 ;
        RECT  6.420 3.440 8.735 3.940 ;
        RECT  6.160 3.285 6.420 3.940 ;
        RECT  3.155 3.440 6.160 3.940 ;
        RECT  2.895 3.285 3.155 3.940 ;
        RECT  0.925 3.440 2.895 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.045 1.565 9.145 1.825 ;
        RECT  8.885 1.565 9.045 2.690 ;
        RECT  7.330 2.530 8.885 2.690 ;
        RECT  7.825 2.870 8.085 3.130 ;
        RECT  7.820 1.035 7.940 1.295 ;
        RECT  7.820 2.090 7.870 2.350 ;
        RECT  6.760 2.870 7.825 3.030 ;
        RECT  7.660 0.615 7.820 2.350 ;
        RECT  6.130 0.615 7.660 0.775 ;
        RECT  7.610 2.090 7.660 2.350 ;
        RECT  7.330 1.035 7.430 1.295 ;
        RECT  7.170 1.035 7.330 2.690 ;
        RECT  7.160 2.280 7.170 2.690 ;
        RECT  7.070 2.280 7.160 2.540 ;
        RECT  6.720 1.035 6.920 1.295 ;
        RECT  6.720 2.125 6.820 2.385 ;
        RECT  6.600 2.735 6.760 3.030 ;
        RECT  6.560 0.955 6.720 2.385 ;
        RECT  5.450 2.735 6.600 2.895 ;
        RECT  5.790 0.955 6.560 1.115 ;
        RECT  5.970 0.530 6.130 0.775 ;
        RECT  4.050 0.530 5.970 0.690 ;
        RECT  5.790 1.295 5.920 1.455 ;
        RECT  5.630 0.885 5.790 1.115 ;
        RECT  5.630 1.295 5.790 2.545 ;
        RECT  4.480 0.885 5.630 1.045 ;
        RECT  5.290 1.275 5.450 2.895 ;
        RECT  5.120 1.275 5.290 1.435 ;
        RECT  4.810 2.735 5.290 2.895 ;
        RECT  4.950 1.615 5.110 2.555 ;
        RECT  4.820 1.615 4.950 1.775 ;
        RECT  4.560 2.395 4.950 2.555 ;
        RECT  4.660 1.225 4.820 1.775 ;
        RECT  4.610 1.955 4.770 2.215 ;
        RECT  4.480 1.955 4.610 2.165 ;
        RECT  4.460 2.395 4.560 2.795 ;
        RECT  4.320 0.885 4.480 2.165 ;
        RECT  4.400 2.395 4.460 3.010 ;
        RECT  4.300 2.535 4.400 3.010 ;
        RECT  4.050 2.005 4.320 2.165 ;
        RECT  2.320 2.850 4.300 3.010 ;
        RECT  3.540 1.485 4.140 1.745 ;
        RECT  3.890 0.530 4.050 1.305 ;
        RECT  3.950 2.005 4.050 2.425 ;
        RECT  3.840 2.005 3.950 2.670 ;
        RECT  3.790 0.755 3.890 1.305 ;
        RECT  3.790 2.165 3.840 2.670 ;
        RECT  2.530 0.755 3.790 0.915 ;
        RECT  2.320 2.510 3.790 2.670 ;
        RECT  3.380 1.095 3.540 2.330 ;
        RECT  2.305 1.095 3.380 1.255 ;
        RECT  2.660 2.170 3.380 2.330 ;
        RECT  2.500 2.015 2.660 2.330 ;
        RECT  2.370 0.695 2.530 0.915 ;
        RECT  2.355 2.015 2.500 2.175 ;
        RECT  1.665 0.695 2.370 0.855 ;
        RECT  2.175 2.380 2.320 2.670 ;
        RECT  2.160 2.850 2.320 3.260 ;
        RECT  2.160 1.595 2.175 2.670 ;
        RECT  2.015 1.595 2.160 2.540 ;
        RECT  1.495 3.100 2.160 3.260 ;
        RECT  2.005 1.595 2.015 1.755 ;
        RECT  1.845 1.045 2.005 1.755 ;
        RECT  1.835 2.760 1.980 2.920 ;
        RECT  1.665 1.965 1.835 2.225 ;
        RECT  1.675 2.480 1.835 2.920 ;
        RECT  1.325 2.480 1.675 2.640 ;
        RECT  1.505 0.695 1.665 2.225 ;
        RECT  1.335 2.945 1.495 3.260 ;
        RECT  0.385 2.945 1.335 3.105 ;
        RECT  1.165 1.035 1.325 2.640 ;
        RECT  1.075 1.035 1.165 1.295 ;
        RECT  1.065 2.070 1.165 2.330 ;
        RECT  0.745 1.500 0.985 1.760 ;
        RECT  0.585 1.135 0.745 2.330 ;
        RECT  0.385 1.135 0.585 1.295 ;
        RECT  0.385 2.170 0.585 2.330 ;
        RECT  0.125 0.695 0.385 1.295 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END ADDFX2

MACRO ADDFX1
    CLASS CORE ;
    FOREIGN ADDFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.325 0.975 9.535 2.375 ;
        RECT  9.275 0.975 9.325 1.235 ;
        RECT  9.275 2.115 9.325 2.375 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.455 1.515 8.615 1.990 ;
        RECT  8.295 0.975 8.455 2.265 ;
        RECT  8.190 0.975 8.295 1.235 ;
        RECT  8.195 2.005 8.295 2.265 ;
        END
        ANTENNADIFFAREA     0.3625 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 2.260 6.320 2.520 ;
        RECT  6.265 1.700 6.315 2.520 ;
        RECT  6.105 1.310 6.265 2.520 ;
        RECT  6.100 1.310 6.105 1.925 ;
        RECT  6.060 2.260 6.105 2.520 ;
        END
        ANTENNAGATEAREA     0.1976 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.490 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.510 3.165 1.990 ;
        RECT  2.645 1.510 2.885 1.825 ;
        END
        ANTENNAGATEAREA     0.2769 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.995 -0.250 9.660 0.250 ;
        RECT  8.735 -0.250 8.995 1.145 ;
        RECT  6.570 -0.250 8.735 0.250 ;
        RECT  6.310 -0.250 6.570 0.405 ;
        RECT  3.115 -0.250 6.310 0.250 ;
        RECT  2.855 -0.250 3.115 0.575 ;
        RECT  0.925 -0.250 2.855 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.995 3.440 9.660 3.940 ;
        RECT  8.735 2.880 8.995 3.940 ;
        RECT  6.420 3.440 8.735 3.940 ;
        RECT  6.160 3.285 6.420 3.940 ;
        RECT  3.155 3.440 6.160 3.940 ;
        RECT  2.895 3.285 3.155 3.940 ;
        RECT  0.925 3.440 2.895 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.045 1.565 9.145 1.825 ;
        RECT  8.885 1.565 9.045 2.690 ;
        RECT  7.330 2.530 8.885 2.690 ;
        RECT  7.825 2.870 8.085 3.130 ;
        RECT  7.820 1.035 7.940 1.295 ;
        RECT  7.820 2.090 7.870 2.350 ;
        RECT  6.760 2.870 7.825 3.030 ;
        RECT  7.660 0.615 7.820 2.350 ;
        RECT  6.130 0.615 7.660 0.775 ;
        RECT  7.610 2.090 7.660 2.350 ;
        RECT  7.330 1.035 7.430 1.295 ;
        RECT  7.170 1.035 7.330 2.690 ;
        RECT  7.160 2.280 7.170 2.690 ;
        RECT  7.070 2.280 7.160 2.540 ;
        RECT  6.720 1.035 6.920 1.295 ;
        RECT  6.720 2.125 6.820 2.385 ;
        RECT  6.600 2.735 6.760 3.030 ;
        RECT  6.560 0.955 6.720 2.385 ;
        RECT  5.450 2.735 6.600 2.895 ;
        RECT  5.790 0.955 6.560 1.115 ;
        RECT  5.970 0.530 6.130 0.775 ;
        RECT  4.050 0.530 5.970 0.690 ;
        RECT  5.790 1.295 5.920 1.455 ;
        RECT  5.630 0.885 5.790 1.115 ;
        RECT  5.630 1.295 5.790 2.545 ;
        RECT  4.480 0.885 5.630 1.045 ;
        RECT  5.290 1.275 5.450 2.895 ;
        RECT  5.120 1.275 5.290 1.435 ;
        RECT  4.810 2.735 5.290 2.895 ;
        RECT  4.950 1.615 5.110 2.555 ;
        RECT  4.820 1.615 4.950 1.775 ;
        RECT  4.560 2.395 4.950 2.555 ;
        RECT  4.660 1.225 4.820 1.775 ;
        RECT  4.480 1.955 4.770 2.215 ;
        RECT  4.460 2.395 4.560 2.795 ;
        RECT  4.320 0.885 4.480 2.215 ;
        RECT  4.400 2.395 4.460 3.010 ;
        RECT  4.300 2.535 4.400 3.010 ;
        RECT  4.050 2.055 4.320 2.215 ;
        RECT  2.320 2.850 4.300 3.010 ;
        RECT  3.540 1.485 4.140 1.745 ;
        RECT  3.890 0.530 4.050 1.305 ;
        RECT  3.950 2.055 4.050 2.425 ;
        RECT  3.840 2.055 3.950 2.670 ;
        RECT  3.790 0.755 3.890 1.305 ;
        RECT  3.790 2.165 3.840 2.670 ;
        RECT  2.530 0.755 3.790 0.915 ;
        RECT  2.320 2.510 3.790 2.670 ;
        RECT  3.380 1.095 3.540 2.330 ;
        RECT  2.305 1.095 3.380 1.255 ;
        RECT  2.660 2.170 3.380 2.330 ;
        RECT  2.500 2.015 2.660 2.330 ;
        RECT  2.370 0.695 2.530 0.915 ;
        RECT  2.355 2.015 2.500 2.175 ;
        RECT  1.665 0.695 2.370 0.855 ;
        RECT  2.175 2.380 2.320 2.670 ;
        RECT  2.160 2.850 2.320 3.260 ;
        RECT  2.160 1.595 2.175 2.670 ;
        RECT  2.015 1.595 2.160 2.540 ;
        RECT  1.495 3.100 2.160 3.260 ;
        RECT  2.005 1.595 2.015 1.755 ;
        RECT  1.845 1.045 2.005 1.755 ;
        RECT  1.835 2.760 1.980 2.920 ;
        RECT  1.665 1.965 1.835 2.225 ;
        RECT  1.675 2.480 1.835 2.920 ;
        RECT  1.325 2.480 1.675 2.640 ;
        RECT  1.505 0.695 1.665 2.225 ;
        RECT  1.335 2.945 1.495 3.260 ;
        RECT  0.385 2.945 1.335 3.105 ;
        RECT  1.165 1.035 1.325 2.640 ;
        RECT  1.075 1.035 1.165 1.295 ;
        RECT  1.065 2.070 1.165 2.640 ;
        RECT  0.745 1.500 0.985 1.760 ;
        RECT  0.585 1.135 0.745 2.330 ;
        RECT  0.385 1.135 0.585 1.295 ;
        RECT  0.385 2.170 0.585 2.330 ;
        RECT  0.125 0.695 0.385 1.295 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END ADDFX1

MACRO ADDFXL
    CLASS CORE ;
    FOREIGN ADDFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.865 1.035 9.075 2.265 ;
        RECT  8.810 1.035 8.865 1.295 ;
        RECT  8.815 2.005 8.865 2.265 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.105 0.620 8.230 1.990 ;
        RECT  8.070 0.620 8.105 2.285 ;
        RECT  8.010 0.620 8.070 0.780 ;
        RECT  7.945 1.700 8.070 2.285 ;
        RECT  7.850 0.515 8.010 0.780 ;
        RECT  7.890 2.025 7.945 2.285 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.310 1.700 6.315 1.990 ;
        RECT  6.210 1.310 6.310 1.990 ;
        RECT  6.105 1.310 6.210 2.520 ;
        RECT  6.050 1.765 6.105 2.520 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.490 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.840 1.635 3.095 1.990 ;
        RECT  2.645 1.635 2.840 1.825 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.670 -0.250 9.200 0.250 ;
        RECT  8.410 -0.250 8.670 0.745 ;
        RECT  6.510 -0.250 8.410 0.250 ;
        RECT  6.250 -0.250 6.510 0.405 ;
        RECT  3.295 -0.250 6.250 0.250 ;
        RECT  3.035 -0.250 3.295 0.575 ;
        RECT  0.785 -0.250 3.035 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.525 3.440 9.200 3.940 ;
        RECT  8.265 2.895 8.525 3.940 ;
        RECT  6.350 3.440 8.265 3.940 ;
        RECT  6.090 3.075 6.350 3.940 ;
        RECT  3.155 3.440 6.090 3.940 ;
        RECT  2.895 3.285 3.155 3.940 ;
        RECT  0.785 3.440 2.895 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.645 2.445 8.905 2.705 ;
        RECT  7.170 2.530 8.645 2.690 ;
        RECT  7.825 2.870 8.085 3.220 ;
        RECT  7.670 1.065 7.890 1.325 ;
        RECT  6.690 3.060 7.825 3.220 ;
        RECT  7.510 0.615 7.670 2.350 ;
        RECT  6.080 0.615 7.510 0.775 ;
        RECT  7.310 2.090 7.510 2.350 ;
        RECT  7.170 1.065 7.330 1.665 ;
        RECT  7.080 1.505 7.170 1.665 ;
        RECT  7.080 2.530 7.170 2.880 ;
        RECT  6.920 1.505 7.080 2.880 ;
        RECT  6.910 2.720 6.920 2.880 ;
        RECT  6.770 1.065 6.870 1.325 ;
        RECT  6.665 0.955 6.770 1.325 ;
        RECT  6.530 2.735 6.690 3.220 ;
        RECT  6.505 0.955 6.665 2.430 ;
        RECT  5.390 2.735 6.530 2.895 ;
        RECT  5.740 0.955 6.505 1.115 ;
        RECT  6.420 2.170 6.505 2.430 ;
        RECT  5.920 0.530 6.080 0.775 ;
        RECT  3.985 0.530 5.920 0.690 ;
        RECT  5.730 1.295 5.920 1.455 ;
        RECT  5.580 0.885 5.740 1.115 ;
        RECT  5.570 1.295 5.730 2.545 ;
        RECT  4.480 0.885 5.580 1.045 ;
        RECT  5.230 1.275 5.390 2.895 ;
        RECT  5.120 1.275 5.230 1.435 ;
        RECT  4.840 2.735 5.230 2.895 ;
        RECT  4.890 1.615 5.050 2.555 ;
        RECT  4.820 1.615 4.890 1.775 ;
        RECT  4.590 2.395 4.890 2.555 ;
        RECT  4.660 1.225 4.820 1.775 ;
        RECT  4.480 1.955 4.710 2.215 ;
        RECT  4.490 2.395 4.590 2.865 ;
        RECT  4.430 2.395 4.490 3.075 ;
        RECT  4.320 0.885 4.480 2.215 ;
        RECT  4.330 2.605 4.430 3.075 ;
        RECT  2.345 2.915 4.330 3.075 ;
        RECT  4.080 2.055 4.320 2.215 ;
        RECT  3.540 1.485 4.140 1.745 ;
        RECT  3.820 2.055 4.080 2.735 ;
        RECT  3.825 0.530 3.985 1.305 ;
        RECT  3.725 0.755 3.825 1.305 ;
        RECT  3.790 2.055 3.820 2.670 ;
        RECT  2.320 2.510 3.790 2.670 ;
        RECT  2.855 0.755 3.725 0.915 ;
        RECT  3.475 1.485 3.540 2.330 ;
        RECT  3.315 1.095 3.475 2.330 ;
        RECT  3.215 1.095 3.315 1.455 ;
        RECT  2.660 2.170 3.315 2.330 ;
        RECT  2.515 1.295 3.215 1.455 ;
        RECT  2.695 0.695 2.855 0.915 ;
        RECT  1.665 0.695 2.695 0.855 ;
        RECT  2.500 2.015 2.660 2.330 ;
        RECT  2.355 1.035 2.515 1.455 ;
        RECT  2.355 2.015 2.500 2.175 ;
        RECT  2.185 2.915 2.345 3.220 ;
        RECT  2.175 2.355 2.320 2.670 ;
        RECT  1.485 3.060 2.185 3.220 ;
        RECT  2.160 1.135 2.175 2.670 ;
        RECT  2.015 1.135 2.160 2.515 ;
        RECT  2.005 1.135 2.015 1.295 ;
        RECT  1.845 1.035 2.005 1.295 ;
        RECT  1.835 2.720 1.980 2.880 ;
        RECT  1.665 1.965 1.835 2.225 ;
        RECT  1.675 2.480 1.835 2.880 ;
        RECT  1.325 2.480 1.675 2.640 ;
        RECT  1.505 0.695 1.665 2.225 ;
        RECT  1.325 2.820 1.485 3.220 ;
        RECT  1.165 1.035 1.325 2.640 ;
        RECT  0.745 2.820 1.325 2.980 ;
        RECT  1.075 1.035 1.165 1.295 ;
        RECT  1.065 2.070 1.165 2.330 ;
        RECT  0.745 1.500 0.985 1.760 ;
        RECT  0.585 1.135 0.745 2.980 ;
        RECT  0.385 1.135 0.585 1.295 ;
        RECT  0.125 2.170 0.585 2.430 ;
        RECT  0.125 1.035 0.385 1.295 ;
    END
END ADDFXL

MACRO ADDHX4
    CLASS CORE ;
    FOREIGN ADDHX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.800 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.130 0.495 8.550 0.800 ;
        RECT  7.530 0.600 8.130 0.800 ;
        RECT  7.590 1.965 7.850 2.225 ;
        RECT  6.830 1.965 7.590 2.165 ;
        RECT  7.270 0.600 7.530 0.890 ;
        RECT  6.510 0.600 7.270 0.800 ;
        RECT  6.775 1.965 6.830 2.565 ;
        RECT  6.570 1.965 6.775 2.810 ;
        RECT  6.565 2.110 6.570 2.810 ;
        RECT  3.145 2.170 6.565 2.370 ;
        RECT  6.250 0.600 6.510 1.300 ;
        RECT  5.490 1.100 6.250 1.300 ;
        RECT  5.230 1.035 5.490 1.300 ;
        RECT  4.485 1.100 5.230 1.300 ;
        RECT  4.365 1.065 4.485 1.300 ;
        RECT  4.205 1.065 4.365 1.445 ;
        RECT  3.145 1.285 4.205 1.445 ;
        RECT  2.985 1.285 3.145 2.370 ;
        END
        ANTENNADIFFAREA     3.7667 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.665 1.515 13.675 2.400 ;
        RECT  13.465 0.915 13.665 2.650 ;
        RECT  13.215 0.915 13.465 1.115 ;
        RECT  13.155 2.450 13.465 2.650 ;
        RECT  13.165 0.695 13.215 1.115 ;
        RECT  12.905 0.495 13.165 1.115 ;
        RECT  12.895 2.450 13.155 3.050 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.735 1.430 7.995 1.785 ;
        RECT  3.555 1.625 7.735 1.785 ;
        RECT  3.345 1.625 3.555 1.990 ;
        RECT  3.325 1.625 3.345 1.785 ;
        END
        ANTENNAGATEAREA     1.7394 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.535 1.620 11.300 1.780 ;
        RECT  9.340 1.290 9.535 1.780 ;
        RECT  9.325 1.290 9.340 1.620 ;
        END
        ANTENNAGATEAREA     1.6705 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.675 -0.250 13.800 0.250 ;
        RECT  13.415 -0.250 13.675 0.705 ;
        RECT  12.655 -0.250 13.415 0.250 ;
        RECT  12.395 -0.250 12.655 0.755 ;
        RECT  11.745 -0.250 12.395 0.250 ;
        RECT  11.485 -0.250 11.745 1.075 ;
        RECT  10.725 -0.250 11.485 0.250 ;
        RECT  10.465 -0.250 10.725 1.075 ;
        RECT  9.810 -0.250 10.465 0.250 ;
        RECT  9.550 -0.250 9.810 0.405 ;
        RECT  3.725 -0.250 9.550 0.250 ;
        RECT  3.465 -0.250 3.725 0.405 ;
        RECT  2.465 -0.250 3.465 0.250 ;
        RECT  2.205 -0.250 2.465 0.405 ;
        RECT  1.405 -0.250 2.205 0.250 ;
        RECT  1.145 -0.250 1.405 0.755 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.665 3.440 13.800 3.940 ;
        RECT  13.405 2.935 13.665 3.940 ;
        RECT  12.645 3.440 13.405 3.940 ;
        RECT  12.385 2.535 12.645 3.940 ;
        RECT  11.625 3.440 12.385 3.940 ;
        RECT  11.365 2.835 11.625 3.940 ;
        RECT  10.570 3.440 11.365 3.940 ;
        RECT  10.310 3.285 10.570 3.940 ;
        RECT  9.470 3.440 10.310 3.940 ;
        RECT  9.210 3.285 9.470 3.940 ;
        RECT  8.415 3.440 9.210 3.940 ;
        RECT  8.155 3.285 8.415 3.940 ;
        RECT  3.255 3.440 8.155 3.940 ;
        RECT  2.995 3.285 3.255 3.940 ;
        RECT  2.455 3.440 2.995 3.940 ;
        RECT  2.195 3.285 2.455 3.940 ;
        RECT  1.405 3.440 2.195 3.940 ;
        RECT  1.145 2.510 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 1.955 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.990 1.295 13.150 2.240 ;
        RECT  12.255 1.295 12.990 1.455 ;
        RECT  12.135 2.080 12.990 2.240 ;
        RECT  11.795 1.635 12.810 1.795 ;
        RECT  12.045 1.035 12.255 1.455 ;
        RECT  11.975 2.080 12.135 3.005 ;
        RECT  11.995 1.035 12.045 1.415 ;
        RECT  11.235 1.255 11.995 1.415 ;
        RECT  11.875 2.405 11.975 3.005 ;
        RECT  11.115 2.405 11.875 2.565 ;
        RECT  11.635 1.635 11.795 2.125 ;
        RECT  8.920 1.965 11.635 2.125 ;
        RECT  10.975 0.610 11.235 1.415 ;
        RECT  10.855 2.405 11.115 3.005 ;
        RECT  10.215 1.255 10.975 1.415 ;
        RECT  10.020 2.405 10.855 2.565 ;
        RECT  10.055 0.865 10.215 1.415 ;
        RECT  9.955 0.865 10.055 1.125 ;
        RECT  9.760 2.310 10.020 2.910 ;
        RECT  8.385 2.750 9.760 2.910 ;
        RECT  8.900 1.035 8.950 1.295 ;
        RECT  8.900 1.965 8.920 2.565 ;
        RECT  8.740 1.035 8.900 2.565 ;
        RECT  8.690 1.035 8.740 1.295 ;
        RECT  8.660 1.965 8.740 2.565 ;
        RECT  8.225 1.075 8.385 2.910 ;
        RECT  8.040 1.075 8.225 1.240 ;
        RECT  7.340 2.595 8.225 2.755 ;
        RECT  7.780 0.980 8.040 1.240 ;
        RECT  7.020 1.080 7.780 1.240 ;
        RECT  7.080 2.595 7.340 3.195 ;
        RECT  6.315 3.035 7.080 3.195 ;
        RECT  6.760 0.980 7.020 1.240 ;
        RECT  6.215 2.935 6.315 3.195 ;
        RECT  6.055 2.605 6.215 3.195 ;
        RECT  2.385 2.605 6.055 2.765 ;
        RECT  5.740 0.495 6.000 0.755 ;
        RECT  4.980 0.535 5.740 0.695 ;
        RECT  1.915 2.945 5.295 3.105 ;
        RECT  4.720 0.495 4.980 0.755 ;
        RECT  1.915 0.585 4.720 0.745 ;
        RECT  2.805 0.925 4.020 1.085 ;
        RECT  2.645 0.925 2.805 2.355 ;
        RECT  2.225 1.685 2.385 2.765 ;
        RECT  2.045 1.685 2.225 1.845 ;
        RECT  1.105 1.585 2.045 1.845 ;
        RECT  1.655 0.585 1.915 1.295 ;
        RECT  1.655 2.165 1.915 3.105 ;
        RECT  0.895 1.135 1.655 1.295 ;
        RECT  0.895 2.165 1.655 2.325 ;
        RECT  0.850 0.695 0.895 1.295 ;
        RECT  0.850 2.165 0.895 3.105 ;
        RECT  0.690 0.695 0.850 3.105 ;
        RECT  0.635 0.695 0.690 1.295 ;
        RECT  0.635 2.165 0.690 3.105 ;
    END
END ADDHX4

MACRO ADDHX2
    CLASS CORE ;
    FOREIGN ADDHX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.425 1.030 4.585 1.290 ;
        RECT  3.615 1.030 4.425 1.190 ;
        RECT  4.135 2.185 4.395 2.445 ;
        RECT  3.990 2.185 4.135 2.400 ;
        RECT  3.555 2.240 3.990 2.400 ;
        RECT  3.355 0.520 3.615 1.190 ;
        RECT  3.375 2.110 3.555 2.400 ;
        RECT  3.345 2.110 3.375 2.715 ;
        RECT  3.345 0.695 3.355 1.190 ;
        RECT  2.595 1.030 3.345 1.190 ;
        RECT  3.115 2.115 3.345 2.715 ;
        RECT  3.070 2.115 3.115 2.400 ;
        RECT  2.495 2.240 3.070 2.400 ;
        RECT  2.495 0.905 2.595 1.190 ;
        RECT  2.335 0.905 2.495 2.400 ;
        RECT  2.095 2.140 2.335 2.400 ;
        END
        ANTENNADIFFAREA     2.1949 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.565 1.105 8.615 2.995 ;
        RECT  8.515 1.105 8.565 3.115 ;
        RECT  8.355 0.645 8.515 3.115 ;
        RECT  8.255 0.645 8.355 1.245 ;
        RECT  8.305 2.175 8.355 3.115 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.470 4.485 1.730 ;
        RECT  4.265 1.470 4.475 1.990 ;
        RECT  4.255 1.470 4.265 1.855 ;
        RECT  3.035 1.695 4.255 1.855 ;
        RECT  2.775 1.595 3.035 1.855 ;
        END
        ANTENNAGATEAREA     0.8853 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.525 7.265 1.785 ;
        RECT  5.670 1.290 5.855 1.785 ;
        RECT  5.645 1.290 5.670 1.580 ;
        END
        ANTENNAGATEAREA     0.8853 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.005 -0.250 8.740 0.250 ;
        RECT  7.745 -0.250 8.005 0.755 ;
        RECT  7.090 -0.250 7.745 0.250 ;
        RECT  6.830 -0.250 7.090 0.815 ;
        RECT  6.030 -0.250 6.830 0.250 ;
        RECT  5.770 -0.250 6.030 0.405 ;
        RECT  1.355 -0.250 5.770 0.250 ;
        RECT  1.195 -0.250 1.355 0.755 ;
        RECT  0.385 -0.250 1.195 0.250 ;
        RECT  0.125 -0.250 0.385 1.095 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.050 3.440 8.740 3.940 ;
        RECT  7.790 2.595 8.050 3.940 ;
        RECT  7.025 3.440 7.790 3.940 ;
        RECT  6.765 2.835 7.025 3.940 ;
        RECT  5.965 3.440 6.765 3.940 ;
        RECT  5.705 3.285 5.965 3.940 ;
        RECT  4.905 3.440 5.705 3.940 ;
        RECT  4.645 3.285 4.905 3.940 ;
        RECT  1.445 3.440 4.645 3.940 ;
        RECT  1.185 3.285 1.445 3.940 ;
        RECT  0.385 3.440 1.185 3.940 ;
        RECT  0.125 2.935 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.940 1.585 8.090 1.845 ;
        RECT  7.780 1.585 7.940 2.170 ;
        RECT  5.460 2.010 7.780 2.170 ;
        RECT  7.340 1.035 7.600 1.295 ;
        RECT  7.275 2.395 7.535 2.995 ;
        RECT  6.580 1.035 7.340 1.220 ;
        RECT  6.515 2.395 7.275 2.555 ;
        RECT  6.320 0.620 6.580 1.220 ;
        RECT  6.255 2.395 6.515 3.095 ;
        RECT  5.610 0.620 6.320 0.780 ;
        RECT  4.925 2.935 6.255 3.095 ;
        RECT  5.450 0.525 5.610 0.780 ;
        RECT  5.270 2.010 5.460 2.565 ;
        RECT  4.925 0.525 5.450 0.685 ;
        RECT  5.200 0.865 5.270 2.565 ;
        RECT  5.110 0.865 5.200 2.170 ;
        RECT  4.765 0.525 4.925 3.095 ;
        RECT  4.125 0.525 4.765 0.685 ;
        RECT  3.885 2.935 4.765 3.095 ;
        RECT  3.865 0.525 4.125 0.785 ;
        RECT  3.625 2.610 3.885 3.210 ;
        RECT  0.915 2.935 3.625 3.095 ;
        RECT  2.845 0.505 3.105 0.795 ;
        RECT  1.405 2.580 2.865 2.740 ;
        RECT  1.695 0.505 2.845 0.665 ;
        RECT  1.875 0.845 2.035 1.635 ;
        RECT  1.845 1.475 1.875 1.635 ;
        RECT  1.685 1.475 1.845 2.215 ;
        RECT  1.535 0.505 1.695 1.290 ;
        RECT  1.585 1.955 1.685 2.215 ;
        RECT  1.405 1.130 1.535 1.290 ;
        RECT  1.245 1.130 1.405 2.740 ;
        RECT  0.895 1.130 1.245 1.290 ;
        RECT  0.635 2.115 1.245 2.375 ;
        RECT  0.450 1.585 1.065 1.845 ;
        RECT  0.755 2.590 0.915 3.095 ;
        RECT  0.635 0.690 0.895 1.290 ;
        RECT  0.450 2.590 0.755 2.750 ;
        RECT  0.290 1.585 0.450 2.750 ;
    END
END ADDHX2

MACRO ADDHX1
    CLASS CORE ;
    FOREIGN ADDHX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.430 1.290 3.555 1.765 ;
        RECT  3.270 1.065 3.430 2.135 ;
        RECT  2.685 1.065 3.270 1.225 ;
        RECT  2.440 1.975 3.270 2.135 ;
        RECT  2.525 0.965 2.685 1.225 ;
        RECT  2.280 1.975 2.440 2.600 ;
        END
        ANTENNADIFFAREA     1.1220 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 1.035 4.990 1.295 ;
        RECT  4.935 1.955 4.990 2.215 ;
        RECT  4.730 1.035 4.935 2.215 ;
        RECT  4.725 1.290 4.730 2.215 ;
        END
        ANTENNADIFFAREA     0.3276 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.110 2.525 4.730 2.685 ;
        RECT  3.950 2.525 4.110 2.940 ;
        RECT  2.100 2.780 3.950 2.940 ;
        RECT  2.930 1.405 3.090 1.795 ;
        RECT  2.100 1.635 2.930 1.795 ;
        RECT  1.940 1.635 2.100 2.940 ;
        RECT  1.715 1.635 1.940 1.795 ;
        RECT  1.505 1.635 1.715 1.990 ;
        RECT  1.285 1.635 1.505 1.895 ;
        END
        ANTENNAGATEAREA     0.4407 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 1.520 4.020 1.990 ;
        END
        ANTENNAGATEAREA     0.4407 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.390 -0.250 5.520 0.250 ;
        RECT  5.130 -0.250 5.390 0.405 ;
        RECT  3.820 -0.250 5.130 0.250 ;
        RECT  3.560 -0.250 3.820 0.405 ;
        RECT  0.925 -0.250 3.560 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.390 3.440 5.520 3.940 ;
        RECT  5.130 3.285 5.390 3.940 ;
        RECT  3.820 3.440 5.130 3.940 ;
        RECT  3.560 3.285 3.820 3.940 ;
        RECT  0.925 3.440 3.560 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.335 1.480 5.375 1.740 ;
        RECT  5.175 0.695 5.335 3.025 ;
        RECT  4.820 0.695 5.175 0.855 ;
        RECT  5.115 1.480 5.175 1.740 ;
        RECT  4.450 2.865 5.175 3.025 ;
        RECT  4.660 0.480 4.820 0.855 ;
        RECT  4.560 0.480 4.660 0.640 ;
        RECT  4.290 2.865 4.450 3.135 ;
        RECT  4.260 1.035 4.360 2.345 ;
        RECT  4.200 0.620 4.260 2.345 ;
        RECT  4.100 0.620 4.200 1.295 ;
        RECT  3.770 2.185 4.200 2.345 ;
        RECT  3.245 0.620 4.100 0.780 ;
        RECT  3.610 2.185 3.770 2.480 ;
        RECT  3.145 2.320 3.610 2.480 ;
        RECT  2.985 0.620 3.245 0.880 ;
        RECT  2.885 2.320 3.145 2.580 ;
        RECT  2.345 0.620 2.985 0.780 ;
        RECT  2.185 0.620 2.345 1.455 ;
        RECT  1.015 1.295 2.185 1.455 ;
        RECT  1.845 0.495 2.005 0.755 ;
        RECT  1.595 0.935 1.855 1.115 ;
        RECT  0.335 0.595 1.845 0.755 ;
        RECT  1.595 2.775 1.755 3.215 ;
        RECT  0.675 0.935 1.595 1.095 ;
        RECT  0.335 2.775 1.595 2.935 ;
        RECT  1.130 2.265 1.390 2.525 ;
        RECT  0.675 2.265 1.130 2.425 ;
        RECT  0.855 1.295 1.015 1.835 ;
        RECT  0.515 0.935 0.675 2.425 ;
        RECT  0.175 0.595 0.335 2.935 ;
    END
END ADDHX1

MACRO ADDHXL
    CLASS CORE ;
    FOREIGN ADDHXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.350 2.110 3.555 2.400 ;
        RECT  3.190 1.915 3.350 2.760 ;
        RECT  3.080 1.915 3.190 2.075 ;
        RECT  2.360 2.600 3.190 2.760 ;
        RECT  2.920 0.575 3.080 2.075 ;
        RECT  1.710 0.575 2.920 0.735 ;
        RECT  2.200 2.210 2.360 2.760 ;
        END
        ANTENNADIFFAREA     0.4379 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.925 0.695 4.935 1.580 ;
        RECT  4.765 0.480 4.925 2.510 ;
        RECT  4.725 0.480 4.765 1.580 ;
        RECT  4.665 2.250 4.765 2.510 ;
        RECT  4.570 0.480 4.725 0.740 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.045 2.650 4.145 2.910 ;
        RECT  3.885 2.650 4.045 3.100 ;
        RECT  2.120 2.940 3.885 3.100 ;
        RECT  2.240 1.260 2.400 2.030 ;
        RECT  2.020 1.870 2.240 2.030 ;
        RECT  2.020 2.940 2.120 3.200 ;
        RECT  1.860 1.870 2.020 3.200 ;
        RECT  1.505 2.110 1.860 2.400 ;
        END
        ANTENNAGATEAREA     0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 1.700 4.015 1.990 ;
        RECT  3.805 1.500 3.965 1.990 ;
        RECT  3.425 1.500 3.805 1.660 ;
        RECT  3.265 1.400 3.425 1.660 ;
        END
        ANTENNAGATEAREA     0.1300 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.255 -0.250 5.060 0.250 ;
        RECT  3.995 -0.250 4.255 0.740 ;
        RECT  3.490 -0.250 3.995 0.250 ;
        RECT  3.230 -0.250 3.490 0.405 ;
        RECT  0.480 -0.250 3.230 0.250 ;
        RECT  0.220 -0.250 0.480 0.405 ;
        RECT  0.000 -0.250 0.220 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.525 3.440 5.060 3.940 ;
        RECT  4.265 3.285 4.525 3.940 ;
        RECT  3.330 3.440 4.265 3.940 ;
        RECT  3.070 3.285 3.330 3.940 ;
        RECT  0.935 3.440 3.070 3.940 ;
        RECT  0.675 3.285 0.935 3.940 ;
        RECT  0.000 3.440 0.675 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.485 1.810 4.575 2.070 ;
        RECT  4.325 1.090 4.485 2.370 ;
        RECT  4.220 1.090 4.325 1.250 ;
        RECT  3.895 2.210 4.325 2.370 ;
        RECT  3.960 0.990 4.220 1.250 ;
        RECT  3.735 2.210 3.895 2.470 ;
        RECT  2.740 2.260 2.930 2.420 ;
        RECT  2.580 0.920 2.740 2.420 ;
        RECT  2.060 0.920 2.580 1.080 ;
        RECT  1.900 0.920 2.060 1.635 ;
        RECT  1.015 1.475 1.900 1.635 ;
        RECT  1.560 0.935 1.720 1.245 ;
        RECT  1.420 2.865 1.680 3.185 ;
        RECT  0.675 1.085 1.560 1.245 ;
        RECT  0.335 2.865 1.420 3.025 ;
        RECT  1.120 0.525 1.380 0.785 ;
        RECT  1.155 2.415 1.315 2.675 ;
        RECT  0.675 2.415 1.155 2.575 ;
        RECT  0.335 0.625 1.120 0.785 ;
        RECT  0.855 1.475 1.015 1.985 ;
        RECT  0.515 1.085 0.675 2.575 ;
        RECT  0.175 0.625 0.335 3.025 ;
    END
END ADDHXL

MACRO TLATNTSCAX20
    CLASS CORE ;
    FOREIGN TLATNTSCAX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.240 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.305 1.765 1.465 ;
        RECT  1.505 1.275 1.715 1.830 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.090 1.105 20.115 2.995 ;
        RECT  19.830 0.720 20.090 3.115 ;
        RECT  19.070 0.720 19.830 2.655 ;
        RECT  18.965 0.720 19.070 3.115 ;
        RECT  16.275 0.720 18.965 1.315 ;
        RECT  18.810 2.045 18.965 3.115 ;
        RECT  18.050 2.045 18.810 2.650 ;
        RECT  17.790 2.045 18.050 3.115 ;
        RECT  17.055 2.045 17.790 2.650 ;
        RECT  16.705 2.045 17.055 3.115 ;
        RECT  16.010 2.045 16.705 2.650 ;
        RECT  11.875 0.715 16.275 1.315 ;
        RECT  15.750 2.045 16.010 3.115 ;
        RECT  15.055 2.045 15.750 2.650 ;
        RECT  14.990 2.045 15.055 2.995 ;
        RECT  14.730 2.045 14.990 3.115 ;
        RECT  13.970 2.045 14.730 2.650 ;
        RECT  13.710 2.045 13.970 3.115 ;
        RECT  12.950 2.045 13.710 2.650 ;
        RECT  12.690 2.045 12.950 3.115 ;
        RECT  11.930 2.045 12.690 2.650 ;
        RECT  11.670 2.045 11.930 3.115 ;
        RECT  11.625 2.335 11.670 2.995 ;
        END
        ANTENNADIFFAREA     5.7648 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 1.700 2.355 1.990 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.575 0.345 2.145 ;
        END
        ANTENNAGATEAREA     0.2574 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.515 -0.250 20.240 0.250 ;
        RECT  11.435 -0.250 19.515 0.405 ;
        RECT  10.825 -0.250 11.435 0.250 ;
        RECT  10.565 -0.250 10.825 0.405 ;
        RECT  9.720 -0.250 10.565 0.250 ;
        RECT  9.460 -0.250 9.720 0.405 ;
        RECT  8.820 -0.250 9.460 0.250 ;
        RECT  8.560 -0.250 8.820 0.405 ;
        RECT  7.665 -0.250 8.560 0.250 ;
        RECT  7.405 -0.250 7.665 0.405 ;
        RECT  6.610 -0.250 7.405 0.250 ;
        RECT  6.010 -0.250 6.610 0.405 ;
        RECT  4.785 -0.250 6.010 0.250 ;
        RECT  4.525 -0.250 4.785 0.405 ;
        RECT  2.895 -0.250 4.525 0.250 ;
        RECT  2.295 -0.250 2.895 0.405 ;
        RECT  1.300 -0.250 2.295 0.250 ;
        RECT  0.700 -0.250 1.300 0.405 ;
        RECT  0.000 -0.250 0.700 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.580 3.440 20.240 3.940 ;
        RECT  19.320 2.895 19.580 3.940 ;
        RECT  18.560 3.440 19.320 3.940 ;
        RECT  18.300 2.895 18.560 3.940 ;
        RECT  17.540 3.440 18.300 3.940 ;
        RECT  17.280 2.895 17.540 3.940 ;
        RECT  16.520 3.440 17.280 3.940 ;
        RECT  16.260 2.895 16.520 3.940 ;
        RECT  15.500 3.440 16.260 3.940 ;
        RECT  15.240 2.895 15.500 3.940 ;
        RECT  14.480 3.440 15.240 3.940 ;
        RECT  14.220 2.895 14.480 3.940 ;
        RECT  13.460 3.440 14.220 3.940 ;
        RECT  13.200 2.895 13.460 3.940 ;
        RECT  12.440 3.440 13.200 3.940 ;
        RECT  12.180 2.895 12.440 3.940 ;
        RECT  11.420 3.440 12.180 3.940 ;
        RECT  11.160 2.255 11.420 3.940 ;
        RECT  10.400 3.440 11.160 3.940 ;
        RECT  10.140 2.255 10.400 3.940 ;
        RECT  9.380 3.440 10.140 3.940 ;
        RECT  9.120 2.425 9.380 3.940 ;
        RECT  8.305 3.440 9.120 3.940 ;
        RECT  8.045 2.400 8.305 3.940 ;
        RECT  6.580 3.440 8.045 3.940 ;
        RECT  6.320 3.285 6.580 3.940 ;
        RECT  5.285 3.440 6.320 3.940 ;
        RECT  5.025 3.390 5.285 3.940 ;
        RECT  4.775 3.440 5.025 3.940 ;
        RECT  4.515 3.285 4.775 3.940 ;
        RECT  3.025 3.440 4.515 3.940 ;
        RECT  2.765 3.285 3.025 3.940 ;
        RECT  1.365 3.440 2.765 3.940 ;
        RECT  1.205 2.905 1.365 3.940 ;
        RECT  0.385 3.440 1.205 3.940 ;
        RECT  0.125 2.845 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.720 1.555 18.460 1.785 ;
        RECT  11.265 1.555 11.720 1.715 ;
        RECT  11.265 0.655 11.315 1.185 ;
        RECT  11.175 0.655 11.265 1.715 ;
        RECT  11.015 0.655 11.175 2.070 ;
        RECT  8.995 0.655 11.015 1.185 ;
        RECT  10.910 1.860 11.015 2.070 ;
        RECT  10.650 1.860 10.910 3.025 ;
        RECT  8.730 1.410 10.765 1.670 ;
        RECT  9.890 1.860 10.650 2.070 ;
        RECT  9.730 1.860 9.890 3.135 ;
        RECT  9.630 2.030 9.730 3.135 ;
        RECT  8.870 2.030 9.630 2.245 ;
        RECT  8.710 2.030 8.870 3.050 ;
        RECT  8.570 0.825 8.730 1.850 ;
        RECT  8.610 2.450 8.710 3.050 ;
        RECT  8.270 0.825 8.570 0.985 ;
        RECT  8.410 1.690 8.570 1.850 ;
        RECT  8.250 1.690 8.410 2.210 ;
        RECT  8.130 1.250 8.390 1.510 ;
        RECT  8.010 0.810 8.270 1.070 ;
        RECT  7.480 2.050 8.250 2.210 ;
        RECT  8.065 1.350 8.130 1.510 ;
        RECT  7.905 1.350 8.065 1.870 ;
        RECT  7.240 0.825 8.010 0.985 ;
        RECT  6.780 1.710 7.905 1.870 ;
        RECT  7.375 1.265 7.665 1.530 ;
        RECT  7.320 2.050 7.480 2.995 ;
        RECT  6.785 1.265 7.375 1.425 ;
        RECT  7.220 2.055 7.320 2.995 ;
        RECT  6.980 0.825 7.240 1.085 ;
        RECT  6.625 0.615 6.785 1.425 ;
        RECT  6.620 1.605 6.780 3.105 ;
        RECT  5.675 0.615 6.625 0.775 ;
        RECT  5.555 2.945 6.620 3.105 ;
        RECT  6.280 1.015 6.440 2.075 ;
        RECT  5.885 1.015 6.280 1.175 ;
        RECT  6.125 1.915 6.280 2.075 ;
        RECT  6.075 1.915 6.125 2.215 ;
        RECT  5.675 1.375 6.095 1.715 ;
        RECT  5.865 1.915 6.075 2.590 ;
        RECT  5.740 2.330 5.865 2.590 ;
        RECT  5.515 0.615 5.675 1.715 ;
        RECT  5.395 2.225 5.555 3.105 ;
        RECT  5.145 0.720 5.515 0.880 ;
        RECT  4.910 1.555 5.515 1.715 ;
        RECT  5.105 2.225 5.395 2.385 ;
        RECT  3.460 2.945 5.395 3.105 ;
        RECT  4.535 1.145 5.295 1.305 ;
        RECT  4.910 2.600 5.215 2.760 ;
        RECT  4.885 0.720 5.145 0.920 ;
        RECT  4.750 1.555 4.910 2.760 ;
        RECT  3.650 0.720 4.885 0.880 ;
        RECT  3.915 2.600 4.750 2.760 ;
        RECT  4.375 1.065 4.535 2.050 ;
        RECT  3.470 1.065 4.375 1.225 ;
        RECT  4.035 1.890 4.375 2.050 ;
        RECT  3.695 1.405 4.095 1.565 ;
        RECT  3.875 1.840 4.035 2.100 ;
        RECT  3.655 2.445 3.915 2.760 ;
        RECT  3.535 1.405 3.695 2.135 ;
        RECT  3.460 1.975 3.535 2.135 ;
        RECT  3.310 0.585 3.470 1.225 ;
        RECT  3.300 1.975 3.460 3.105 ;
        RECT  1.325 0.585 3.310 0.745 ;
        RECT  2.530 2.945 3.300 3.105 ;
        RECT  3.100 1.435 3.205 1.695 ;
        RECT  2.940 0.995 3.100 2.720 ;
        RECT  2.315 0.995 2.940 1.155 ;
        RECT  2.155 2.560 2.940 2.720 ;
        RECT  2.585 1.345 2.745 2.340 ;
        RECT  2.535 1.345 2.585 1.670 ;
        RECT  2.135 2.180 2.585 2.340 ;
        RECT  2.120 1.345 2.535 1.505 ;
        RECT  2.370 2.945 2.530 3.260 ;
        RECT  1.705 3.100 2.370 3.260 ;
        RECT  1.995 2.560 2.155 2.920 ;
        RECT  1.960 0.925 2.120 1.505 ;
        RECT  1.895 2.760 1.995 2.920 ;
        RECT  1.685 0.925 1.960 1.085 ;
        RECT  1.545 2.485 1.705 3.260 ;
        RECT  0.895 2.485 1.545 2.645 ;
        RECT  1.165 0.585 1.325 2.115 ;
        RECT  1.045 1.955 1.165 2.115 ;
        RECT  0.885 1.955 1.045 2.215 ;
        RECT  0.765 1.470 0.985 1.750 ;
        RECT  0.695 2.485 0.895 3.160 ;
        RECT  0.695 1.005 0.765 1.750 ;
        RECT  0.635 1.005 0.695 3.160 ;
        RECT  0.605 1.005 0.635 2.645 ;
        RECT  0.385 1.005 0.605 1.165 ;
        RECT  0.535 1.590 0.605 2.645 ;
        RECT  0.125 0.565 0.385 1.165 ;
    END
END TLATNTSCAX20

MACRO TLATNTSCAX16
    CLASS CORE ;
    FOREIGN TLATNTSCAX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.020 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.275 1.745 1.535 ;
        RECT  1.505 1.275 1.715 1.830 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.885 0.880 16.895 2.995 ;
        RECT  16.625 0.710 16.885 3.115 ;
        RECT  16.200 0.710 16.625 2.650 ;
        RECT  15.865 0.705 16.200 2.650 ;
        RECT  15.760 0.705 15.865 3.115 ;
        RECT  9.645 0.705 15.760 1.305 ;
        RECT  15.605 2.045 15.760 3.115 ;
        RECT  14.870 2.045 15.605 2.650 ;
        RECT  14.520 2.045 14.870 3.115 ;
        RECT  13.825 2.045 14.520 2.650 ;
        RECT  13.565 2.045 13.825 3.115 ;
        RECT  12.805 2.045 13.565 2.650 ;
        RECT  12.545 2.045 12.805 3.115 ;
        RECT  11.835 2.045 12.545 2.650 ;
        RECT  11.785 2.045 11.835 2.995 ;
        RECT  11.525 2.045 11.785 3.115 ;
        RECT  10.765 2.045 11.525 2.650 ;
        RECT  10.505 2.045 10.765 3.115 ;
        RECT  9.745 2.045 10.505 2.650 ;
        RECT  9.485 2.045 9.745 3.115 ;
        END
        ANTENNADIFFAREA     5.2008 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 1.825 2.380 2.035 ;
        RECT  2.175 1.755 2.230 2.035 ;
        RECT  1.965 1.700 2.175 2.035 ;
        RECT  1.940 1.825 1.965 2.035 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.765 0.370 2.075 ;
        RECT  0.125 1.575 0.345 2.145 ;
        END
        ANTENNAGATEAREA     0.2145 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.325 -0.250 17.020 0.250 ;
        RECT  9.265 -0.250 16.325 0.405 ;
        RECT  8.505 -0.250 9.265 0.250 ;
        RECT  8.245 -0.250 8.505 0.405 ;
        RECT  7.530 -0.250 8.245 0.250 ;
        RECT  7.270 -0.250 7.530 0.405 ;
        RECT  6.505 -0.250 7.270 0.250 ;
        RECT  6.245 -0.250 6.505 0.405 ;
        RECT  5.450 -0.250 6.245 0.250 ;
        RECT  4.730 -0.250 5.450 0.405 ;
        RECT  2.925 -0.250 4.730 0.250 ;
        RECT  2.325 -0.250 2.925 0.405 ;
        RECT  1.275 -0.250 2.325 0.250 ;
        RECT  0.935 -0.250 1.275 0.405 ;
        RECT  0.675 -0.250 0.935 0.755 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.375 3.440 17.020 3.940 ;
        RECT  16.115 2.895 16.375 3.940 ;
        RECT  15.355 3.440 16.115 3.940 ;
        RECT  15.095 2.895 15.355 3.940 ;
        RECT  14.335 3.440 15.095 3.940 ;
        RECT  14.075 2.895 14.335 3.940 ;
        RECT  13.315 3.440 14.075 3.940 ;
        RECT  13.055 2.895 13.315 3.940 ;
        RECT  12.295 3.440 13.055 3.940 ;
        RECT  12.035 2.895 12.295 3.940 ;
        RECT  11.275 3.440 12.035 3.940 ;
        RECT  11.015 2.895 11.275 3.940 ;
        RECT  10.255 3.440 11.015 3.940 ;
        RECT  9.995 2.895 10.255 3.940 ;
        RECT  9.235 3.440 9.995 3.940 ;
        RECT  8.975 2.595 9.235 3.940 ;
        RECT  8.215 3.440 8.975 3.940 ;
        RECT  7.955 2.595 8.215 3.940 ;
        RECT  7.140 3.440 7.955 3.940 ;
        RECT  6.880 2.400 7.140 3.940 ;
        RECT  5.365 3.440 6.880 3.940 ;
        RECT  5.105 3.285 5.365 3.940 ;
        RECT  3.080 3.440 5.105 3.940 ;
        RECT  2.820 3.285 3.080 3.940 ;
        RECT  1.490 3.440 2.820 3.940 ;
        RECT  1.330 2.905 1.490 3.940 ;
        RECT  0.510 3.440 1.330 3.940 ;
        RECT  0.250 2.845 0.510 3.940 ;
        RECT  0.000 3.440 0.250 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.265 1.615 15.470 1.825 ;
        RECT  9.400 1.555 15.265 1.825 ;
        RECT  9.305 0.680 9.400 1.825 ;
        RECT  9.145 0.680 9.305 2.415 ;
        RECT  7.780 0.680 9.145 1.270 ;
        RECT  8.725 2.075 9.145 2.415 ;
        RECT  7.570 1.510 8.935 1.770 ;
        RECT  8.465 2.075 8.725 3.135 ;
        RECT  7.740 2.075 8.465 2.415 ;
        RECT  7.705 2.075 7.740 2.725 ;
        RECT  7.580 2.075 7.705 3.050 ;
        RECT  7.445 2.450 7.580 3.050 ;
        RECT  7.410 0.905 7.570 1.770 ;
        RECT  7.055 0.905 7.410 1.065 ;
        RECT  7.400 1.610 7.410 1.770 ;
        RECT  7.240 1.610 7.400 2.210 ;
        RECT  6.315 2.050 7.240 2.210 ;
        RECT  7.035 1.265 7.205 1.425 ;
        RECT  6.795 0.805 7.055 1.065 ;
        RECT  6.875 1.265 7.035 1.855 ;
        RECT  5.615 1.695 6.875 1.855 ;
        RECT  6.015 0.905 6.795 1.065 ;
        RECT  6.190 1.310 6.450 1.495 ;
        RECT  6.155 2.050 6.315 2.850 ;
        RECT  5.650 1.310 6.190 1.470 ;
        RECT  6.055 2.250 6.155 2.850 ;
        RECT  5.855 0.870 6.015 1.130 ;
        RECT  5.490 0.600 5.650 1.470 ;
        RECT  5.455 1.655 5.615 3.095 ;
        RECT  4.570 0.600 5.490 0.760 ;
        RECT  4.375 2.935 5.455 3.095 ;
        RECT  5.115 1.070 5.275 2.075 ;
        RECT  4.980 1.070 5.115 1.230 ;
        RECT  4.970 1.915 5.115 2.075 ;
        RECT  4.820 0.965 4.980 1.230 ;
        RECT  4.920 1.915 4.970 2.215 ;
        RECT  4.570 1.455 4.935 1.715 ;
        RECT  4.710 1.915 4.920 2.590 ;
        RECT  4.510 2.310 4.710 2.590 ;
        RECT  4.505 0.600 4.570 1.715 ;
        RECT  4.410 0.600 4.505 2.120 ;
        RECT  3.955 0.660 4.410 0.820 ;
        RECT  4.345 1.505 4.410 2.120 ;
        RECT  4.215 2.935 4.375 3.215 ;
        RECT  3.970 1.960 4.345 2.120 ;
        RECT  3.525 3.055 4.215 3.215 ;
        RECT  3.985 1.030 4.145 1.745 ;
        RECT  3.470 1.030 3.985 1.190 ;
        RECT  3.810 1.960 3.970 2.860 ;
        RECT  3.695 0.560 3.955 0.820 ;
        RECT  3.710 2.260 3.810 2.860 ;
        RECT  3.525 1.405 3.715 1.565 ;
        RECT  3.365 1.405 3.525 3.215 ;
        RECT  3.310 0.585 3.470 1.190 ;
        RECT  2.635 2.935 3.365 3.095 ;
        RECT  1.325 0.585 3.310 0.745 ;
        RECT  3.080 1.665 3.155 1.925 ;
        RECT  2.920 0.995 3.080 2.720 ;
        RECT  2.345 0.995 2.920 1.155 ;
        RECT  2.280 2.560 2.920 2.720 ;
        RECT  2.560 1.345 2.720 2.375 ;
        RECT  2.475 2.935 2.635 3.260 ;
        RECT  2.450 1.345 2.560 1.605 ;
        RECT  2.175 2.215 2.560 2.375 ;
        RECT  1.830 3.100 2.475 3.260 ;
        RECT  2.120 1.345 2.450 1.505 ;
        RECT  2.120 2.560 2.280 2.920 ;
        RECT  1.960 0.925 2.120 1.505 ;
        RECT  2.015 2.760 2.120 2.920 ;
        RECT  1.685 0.925 1.960 1.085 ;
        RECT  1.670 2.485 1.830 3.260 ;
        RECT  1.020 2.485 1.670 2.645 ;
        RECT  1.165 0.585 1.325 2.115 ;
        RECT  1.050 1.955 1.165 2.115 ;
        RECT  0.890 1.955 1.050 2.215 ;
        RECT  0.760 2.485 1.020 3.160 ;
        RECT  0.765 1.490 0.985 1.750 ;
        RECT  0.710 1.130 0.765 1.750 ;
        RECT  0.710 2.485 0.760 2.645 ;
        RECT  0.605 1.130 0.710 2.645 ;
        RECT  0.385 1.130 0.605 1.290 ;
        RECT  0.550 1.590 0.605 2.645 ;
        RECT  0.125 0.690 0.385 1.290 ;
    END
END TLATNTSCAX16

MACRO TLATNTSCAX12
    CLASS CORE ;
    FOREIGN TLATNTSCAX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.275 1.745 1.535 ;
        RECT  1.505 1.275 1.715 1.830 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.995 2.335 14.135 2.585 ;
        RECT  13.795 0.705 14.130 1.305 ;
        RECT  13.990 1.925 13.995 2.650 ;
        RECT  13.795 1.925 13.990 3.115 ;
        RECT  13.640 0.705 13.795 3.115 ;
        RECT  12.965 0.705 13.640 2.650 ;
        RECT  8.530 0.705 12.965 1.305 ;
        RECT  12.945 2.045 12.965 2.650 ;
        RECT  12.685 2.045 12.945 3.115 ;
        RECT  11.925 2.045 12.685 2.650 ;
        RECT  11.665 2.045 11.925 3.115 ;
        RECT  11.625 2.045 11.665 2.995 ;
        RECT  10.915 2.045 11.625 2.650 ;
        RECT  10.905 2.045 10.915 2.995 ;
        RECT  10.645 2.045 10.905 3.115 ;
        RECT  9.885 2.045 10.645 2.650 ;
        RECT  9.625 2.045 9.885 3.115 ;
        RECT  8.865 2.045 9.625 2.650 ;
        RECT  8.605 2.045 8.865 3.115 ;
        END
        ANTENNADIFFAREA     3.9040 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 1.825 2.380 2.035 ;
        RECT  2.175 1.755 2.230 2.035 ;
        RECT  1.965 1.700 2.175 2.035 ;
        RECT  1.940 1.825 1.965 2.035 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.765 0.370 2.045 ;
        RECT  0.125 1.575 0.345 2.145 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.615 -0.250 14.260 0.250 ;
        RECT  13.355 -0.250 13.615 0.405 ;
        RECT  12.585 -0.250 13.355 0.250 ;
        RECT  12.325 -0.250 12.585 0.405 ;
        RECT  11.570 -0.250 12.325 0.250 ;
        RECT  11.310 -0.250 11.570 0.405 ;
        RECT  10.515 -0.250 11.310 0.250 ;
        RECT  10.255 -0.250 10.515 0.405 ;
        RECT  9.480 -0.250 10.255 0.250 ;
        RECT  9.220 -0.250 9.480 0.405 ;
        RECT  8.445 -0.250 9.220 0.250 ;
        RECT  8.185 -0.250 8.445 0.405 ;
        RECT  7.430 -0.250 8.185 0.250 ;
        RECT  7.170 -0.250 7.430 0.405 ;
        RECT  6.385 -0.250 7.170 0.250 ;
        RECT  6.125 -0.250 6.385 0.405 ;
        RECT  5.295 -0.250 6.125 0.250 ;
        RECT  4.575 -0.250 5.295 0.405 ;
        RECT  2.925 -0.250 4.575 0.250 ;
        RECT  2.325 -0.250 2.925 0.405 ;
        RECT  1.275 -0.250 2.325 0.250 ;
        RECT  0.935 -0.250 1.275 0.405 ;
        RECT  0.675 -0.250 0.935 0.755 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.455 3.440 14.260 3.940 ;
        RECT  13.195 2.895 13.455 3.940 ;
        RECT  12.435 3.440 13.195 3.940 ;
        RECT  12.175 2.895 12.435 3.940 ;
        RECT  11.415 3.440 12.175 3.940 ;
        RECT  11.155 2.895 11.415 3.940 ;
        RECT  10.395 3.440 11.155 3.940 ;
        RECT  10.135 2.895 10.395 3.940 ;
        RECT  9.375 3.440 10.135 3.940 ;
        RECT  9.115 2.895 9.375 3.940 ;
        RECT  8.355 3.440 9.115 3.940 ;
        RECT  8.095 2.105 8.355 3.940 ;
        RECT  7.335 3.440 8.095 3.940 ;
        RECT  7.075 2.595 7.335 3.940 ;
        RECT  5.455 3.440 7.075 3.940 ;
        RECT  5.195 3.285 5.455 3.940 ;
        RECT  3.075 3.440 5.195 3.940 ;
        RECT  2.815 3.285 3.075 3.940 ;
        RECT  1.495 3.440 2.815 3.940 ;
        RECT  1.235 2.860 1.495 3.940 ;
        RECT  0.410 3.440 1.235 3.940 ;
        RECT  0.150 2.905 0.410 3.940 ;
        RECT  0.000 3.440 0.150 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.935 1.555 12.455 1.715 ;
        RECT  7.855 0.925 7.935 1.715 ;
        RECT  7.845 0.925 7.855 2.350 ;
        RECT  7.695 0.925 7.845 3.045 ;
        RECT  7.675 0.925 7.695 1.185 ;
        RECT  7.585 2.105 7.695 3.045 ;
        RECT  6.895 1.025 7.675 1.185 ;
        RECT  6.825 2.195 7.585 2.355 ;
        RECT  6.960 1.490 7.430 1.650 ;
        RECT  6.800 1.490 6.960 1.945 ;
        RECT  6.635 0.925 6.895 1.185 ;
        RECT  6.565 2.195 6.825 3.135 ;
        RECT  6.315 1.785 6.800 1.945 ;
        RECT  6.330 1.420 6.380 1.580 ;
        RECT  6.170 0.595 6.330 1.580 ;
        RECT  6.055 1.785 6.315 3.045 ;
        RECT  4.415 0.595 6.170 0.755 ;
        RECT  6.120 1.420 6.170 1.580 ;
        RECT  5.940 1.785 6.055 1.945 ;
        RECT  5.835 1.020 5.940 1.945 ;
        RECT  5.780 0.970 5.835 1.945 ;
        RECT  5.575 0.970 5.780 1.230 ;
        RECT  5.440 1.555 5.600 3.095 ;
        RECT  4.375 2.935 5.440 3.095 ;
        RECT  5.100 1.070 5.260 2.075 ;
        RECT  4.855 1.070 5.100 1.230 ;
        RECT  4.970 1.915 5.100 2.075 ;
        RECT  4.760 1.915 4.970 2.215 ;
        RECT  4.415 1.455 4.920 1.715 ;
        RECT  4.595 0.970 4.855 1.230 ;
        RECT  4.600 1.915 4.760 2.590 ;
        RECT  4.255 0.595 4.415 2.420 ;
        RECT  4.215 2.935 4.375 3.215 ;
        RECT  3.955 0.610 4.255 0.820 ;
        RECT  3.970 2.260 4.255 2.420 ;
        RECT  3.525 3.055 4.215 3.215 ;
        RECT  3.915 1.005 4.075 2.075 ;
        RECT  3.710 2.260 3.970 2.860 ;
        RECT  3.695 0.560 3.955 0.820 ;
        RECT  3.470 1.005 3.915 1.165 ;
        RECT  3.765 1.815 3.915 2.075 ;
        RECT  3.525 1.355 3.730 1.515 ;
        RECT  3.365 1.355 3.525 3.215 ;
        RECT  3.310 0.585 3.470 1.165 ;
        RECT  2.625 2.935 3.365 3.095 ;
        RECT  1.325 0.585 3.310 0.745 ;
        RECT  3.080 1.835 3.180 2.095 ;
        RECT  2.920 1.000 3.080 2.735 ;
        RECT  2.305 1.000 2.920 1.160 ;
        RECT  2.285 2.575 2.920 2.735 ;
        RECT  2.560 1.345 2.720 2.375 ;
        RECT  2.465 2.935 2.625 3.260 ;
        RECT  2.460 1.345 2.560 1.615 ;
        RECT  2.175 2.215 2.560 2.375 ;
        RECT  1.835 3.100 2.465 3.260 ;
        RECT  2.120 1.345 2.460 1.505 ;
        RECT  2.125 2.575 2.285 2.920 ;
        RECT  2.025 2.760 2.125 2.920 ;
        RECT  1.960 0.925 2.120 1.505 ;
        RECT  1.685 0.925 1.960 1.085 ;
        RECT  1.675 2.485 1.835 3.260 ;
        RECT  0.920 2.485 1.675 2.645 ;
        RECT  1.165 0.585 1.325 2.135 ;
        RECT  1.050 1.975 1.165 2.135 ;
        RECT  0.890 1.975 1.050 2.235 ;
        RECT  0.765 1.490 0.985 1.750 ;
        RECT  0.710 2.485 0.920 3.160 ;
        RECT  0.710 1.060 0.765 1.750 ;
        RECT  0.660 1.060 0.710 3.160 ;
        RECT  0.605 1.060 0.660 2.645 ;
        RECT  0.385 1.060 0.605 1.220 ;
        RECT  0.550 1.590 0.605 2.645 ;
        RECT  0.125 0.960 0.385 1.220 ;
    END
END TLATNTSCAX12

MACRO TLATNTSCAX8
    CLASS CORE ;
    FOREIGN TLATNTSCAX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.805 1.425 3.095 1.995 ;
        END
        ANTENNAGATEAREA     0.2002 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.955 0.515 17.355 3.020 ;
        RECT  16.375 0.515 16.955 0.765 ;
        RECT  16.225 2.010 16.955 2.810 ;
        RECT  11.600 0.605 16.375 0.765 ;
        RECT  15.790 2.010 16.225 2.390 ;
        RECT  15.690 2.010 15.790 2.400 ;
        RECT  15.290 2.010 15.690 3.035 ;
        RECT  14.135 2.010 15.290 2.390 ;
        RECT  13.950 2.010 14.135 2.585 ;
        RECT  13.550 2.010 13.950 3.035 ;
        RECT  13.465 2.010 13.550 2.585 ;
        RECT  12.295 2.010 13.465 2.390 ;
        RECT  12.120 2.010 12.295 2.585 ;
        RECT  11.720 2.010 12.120 3.065 ;
        END
        ANTENNADIFFAREA     2.7652 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.370 1.290 3.615 1.940 ;
        RECT  3.345 1.290 3.370 1.720 ;
        END
        ANTENNAGATEAREA     0.2002 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 1.505 1.165 1.765 ;
        RECT  0.795 1.505 0.945 1.925 ;
        RECT  0.585 1.505 0.795 1.990 ;
        RECT  0.565 1.505 0.585 1.765 ;
        END
        ANTENNAGATEAREA     0.8268 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.150 -0.250 17.480 0.250 ;
        RECT  15.890 -0.250 16.150 0.405 ;
        RECT  15.060 -0.250 15.890 0.250 ;
        RECT  14.800 -0.250 15.060 0.405 ;
        RECT  13.860 -0.250 14.800 0.250 ;
        RECT  13.260 -0.250 13.860 0.405 ;
        RECT  12.400 -0.250 13.260 0.250 ;
        RECT  12.140 -0.250 12.400 0.405 ;
        RECT  11.310 -0.250 12.140 0.250 ;
        RECT  11.050 -0.250 11.310 0.405 ;
        RECT  8.830 -0.250 11.050 0.250 ;
        RECT  8.570 -0.250 8.830 0.775 ;
        RECT  7.070 -0.250 8.570 0.250 ;
        RECT  6.810 -0.250 7.070 0.910 ;
        RECT  5.145 -0.250 6.810 0.250 ;
        RECT  4.885 -0.250 5.145 0.405 ;
        RECT  4.045 -0.250 4.885 0.250 ;
        RECT  3.785 -0.250 4.045 0.405 ;
        RECT  2.940 -0.250 3.785 0.250 ;
        RECT  2.680 -0.250 2.940 0.405 ;
        RECT  1.915 -0.250 2.680 0.250 ;
        RECT  1.655 -0.250 1.915 0.910 ;
        RECT  0.895 -0.250 1.655 0.250 ;
        RECT  0.635 -0.250 0.895 1.205 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.480 3.440 17.480 3.940 ;
        RECT  16.220 3.285 16.480 3.940 ;
        RECT  14.770 3.440 16.220 3.940 ;
        RECT  14.510 2.785 14.770 3.940 ;
        RECT  12.990 3.440 14.510 3.940 ;
        RECT  12.730 2.785 12.990 3.940 ;
        RECT  11.095 3.440 12.730 3.940 ;
        RECT  10.835 3.285 11.095 3.940 ;
        RECT  8.965 3.440 10.835 3.940 ;
        RECT  8.705 3.285 8.965 3.940 ;
        RECT  7.195 3.440 8.705 3.940 ;
        RECT  6.935 3.285 7.195 3.940 ;
        RECT  5.210 3.440 6.935 3.940 ;
        RECT  4.950 3.285 5.210 3.940 ;
        RECT  4.110 3.440 4.950 3.940 ;
        RECT  3.850 3.285 4.110 3.940 ;
        RECT  2.880 3.440 3.850 3.940 ;
        RECT  2.620 3.285 2.880 3.940 ;
        RECT  1.955 3.440 2.620 3.940 ;
        RECT  1.695 3.285 1.955 3.940 ;
        RECT  0.895 3.440 1.695 3.940 ;
        RECT  0.635 2.930 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.625 1.260 16.725 1.520 ;
        RECT  16.465 0.945 16.625 1.790 ;
        RECT  11.420 0.945 16.465 1.105 ;
        RECT  11.960 1.630 16.465 1.790 ;
        RECT  11.490 1.290 16.200 1.450 ;
        RECT  11.330 1.290 11.490 2.970 ;
        RECT  11.260 0.630 11.420 1.105 ;
        RECT  10.645 2.810 11.330 2.970 ;
        RECT  10.300 0.630 11.260 0.790 ;
        RECT  10.920 1.045 11.080 2.135 ;
        RECT  10.580 1.045 10.920 1.205 ;
        RECT  10.760 1.975 10.920 2.135 ;
        RECT  10.490 1.975 10.760 2.615 ;
        RECT  10.300 1.475 10.730 1.735 ;
        RECT  10.485 2.810 10.645 3.100 ;
        RECT  10.105 2.940 10.485 3.100 ;
        RECT  10.140 0.630 10.300 2.760 ;
        RECT  9.730 0.630 10.140 0.900 ;
        RECT  5.975 2.600 10.140 2.760 ;
        RECT  9.845 2.940 10.105 3.200 ;
        RECT  9.800 1.435 9.960 2.420 ;
        RECT  5.785 2.940 9.845 3.100 ;
        RECT  9.520 1.435 9.800 1.595 ;
        RECT  5.785 2.260 9.800 2.420 ;
        RECT  9.630 0.630 9.730 1.000 ;
        RECT  9.470 0.630 9.630 1.150 ;
        RECT  9.455 1.810 9.615 2.080 ;
        RECT  9.260 1.335 9.520 1.595 ;
        RECT  7.920 0.990 9.470 1.150 ;
        RECT  8.275 1.810 9.455 1.970 ;
        RECT  7.775 1.355 9.260 1.515 ;
        RECT  8.015 1.710 8.275 1.970 ;
        RECT  5.925 1.810 8.015 1.970 ;
        RECT  7.660 0.870 7.920 1.150 ;
        RECT  7.615 1.355 7.775 1.610 ;
        RECT  7.410 0.990 7.660 1.150 ;
        RECT  6.145 1.450 7.615 1.610 ;
        RECT  7.250 0.990 7.410 1.260 ;
        RECT  6.095 1.100 7.250 1.260 ;
        RECT  5.935 0.705 6.095 1.260 ;
        RECT  5.875 1.710 5.925 1.970 ;
        RECT  5.750 1.710 5.875 2.055 ;
        RECT  5.625 2.260 5.785 3.100 ;
        RECT  5.590 0.930 5.750 2.055 ;
        RECT  1.405 2.940 5.625 3.100 ;
        RECT  5.455 0.930 5.590 1.090 ;
        RECT  5.300 1.895 5.590 2.055 ;
        RECT  5.295 0.585 5.455 1.090 ;
        RECT  4.960 1.400 5.395 1.660 ;
        RECT  5.140 1.895 5.300 2.715 ;
        RECT  2.560 0.585 5.295 0.745 ;
        RECT  2.330 2.555 5.140 2.715 ;
        RECT  4.955 0.990 4.960 1.660 ;
        RECT  4.795 0.990 4.955 2.290 ;
        RECT  4.335 0.990 4.795 1.150 ;
        RECT  4.400 2.130 4.795 2.290 ;
        RECT  4.135 1.620 4.615 1.880 ;
        RECT  3.985 0.930 4.135 1.880 ;
        RECT  3.975 0.930 3.985 2.335 ;
        RECT  3.235 0.930 3.975 1.090 ;
        RECT  3.825 1.720 3.975 2.335 ;
        RECT  3.490 2.175 3.825 2.335 ;
        RECT  2.400 0.585 2.560 2.120 ;
        RECT  2.165 0.695 2.400 1.295 ;
        RECT  2.330 1.960 2.400 2.120 ;
        RECT  2.170 1.960 2.330 2.715 ;
        RECT  2.070 1.960 2.170 2.560 ;
        RECT  1.815 1.480 2.160 1.740 ;
        RECT  1.765 1.480 1.815 2.615 ;
        RECT  1.655 1.150 1.765 2.615 ;
        RECT  1.605 1.150 1.655 1.740 ;
        RECT  1.405 2.455 1.655 2.615 ;
        RECT  1.405 1.150 1.605 1.310 ;
        RECT  1.195 0.615 1.405 1.310 ;
        RECT  1.245 2.065 1.405 3.100 ;
        RECT  1.145 2.065 1.245 3.005 ;
        RECT  1.145 0.615 1.195 1.215 ;
        RECT  0.385 2.455 1.145 2.615 ;
        RECT  0.335 0.620 0.385 1.220 ;
        RECT  0.335 2.065 0.385 3.005 ;
        RECT  0.175 0.620 0.335 3.005 ;
        RECT  0.125 0.620 0.175 1.220 ;
        RECT  0.125 2.065 0.175 3.005 ;
    END
END TLATNTSCAX8

MACRO TLATNTSCAX6
    CLASS CORE ;
    FOREIGN TLATNTSCAX6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.040 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.265 1.295 2.370 1.455 ;
        RECT  2.175 1.295 2.265 1.925 ;
        RECT  2.105 1.295 2.175 1.990 ;
        RECT  1.965 1.700 2.105 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.915 0.585 10.930 2.360 ;
        RECT  10.690 0.585 10.915 2.810 ;
        RECT  8.630 0.585 10.690 0.845 ;
        RECT  10.635 2.110 10.690 2.810 ;
        RECT  10.375 2.110 10.635 3.145 ;
        RECT  10.245 2.110 10.375 2.810 ;
        RECT  9.075 2.115 10.245 2.445 ;
        RECT  8.960 2.115 9.075 2.585 ;
        RECT  8.700 2.115 8.960 3.115 ;
        END
        ANTENNADIFFAREA     1.3520 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.700 2.835 2.270 ;
        RECT  2.595 1.700 2.635 2.400 ;
        RECT  2.425 2.110 2.595 2.400 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 1.575 0.805 2.145 ;
        RECT  0.585 1.470 0.785 2.145 ;
        RECT  0.575 1.470 0.585 1.925 ;
        RECT  0.525 1.470 0.575 1.765 ;
        END
        ANTENNAGATEAREA     0.4251 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.490 -0.250 11.040 0.250 ;
        RECT  10.230 -0.250 10.490 0.405 ;
        RECT  9.390 -0.250 10.230 0.250 ;
        RECT  9.130 -0.250 9.390 0.405 ;
        RECT  8.290 -0.250 9.130 0.250 ;
        RECT  8.030 -0.250 8.290 0.405 ;
        RECT  5.530 -0.250 8.030 0.250 ;
        RECT  5.270 -0.250 5.530 0.405 ;
        RECT  3.155 -0.250 5.270 0.250 ;
        RECT  2.895 -0.250 3.155 0.405 ;
        RECT  1.835 -0.250 2.895 0.250 ;
        RECT  1.235 -0.250 1.835 0.405 ;
        RECT  0.435 -0.250 1.235 0.250 ;
        RECT  0.175 -0.250 0.435 1.280 ;
        RECT  0.000 -0.250 0.175 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.780 3.440 11.040 3.940 ;
        RECT  9.520 2.935 9.780 3.940 ;
        RECT  8.005 3.440 9.520 3.940 ;
        RECT  7.745 2.945 8.005 3.940 ;
        RECT  5.880 3.440 7.745 3.940 ;
        RECT  5.620 3.285 5.880 3.940 ;
        RECT  4.125 3.440 5.620 3.940 ;
        RECT  3.865 3.285 4.125 3.940 ;
        RECT  1.455 3.440 3.865 3.940 ;
        RECT  1.195 2.870 1.455 3.940 ;
        RECT  0.385 3.440 1.195 3.940 ;
        RECT  0.125 2.225 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.425 1.660 10.510 1.920 ;
        RECT  10.350 1.030 10.425 1.920 ;
        RECT  10.265 1.030 10.350 1.880 ;
        RECT  8.450 1.030 10.265 1.190 ;
        RECT  8.770 1.720 10.265 1.880 ;
        RECT  8.430 1.370 10.080 1.530 ;
        RECT  8.290 0.600 8.450 1.190 ;
        RECT  8.270 1.370 8.430 2.745 ;
        RECT  6.935 0.600 8.290 0.760 ;
        RECT  7.455 2.585 8.270 2.745 ;
        RECT  7.930 1.055 8.090 2.135 ;
        RECT  7.290 1.055 7.930 1.215 ;
        RECT  7.670 1.975 7.930 2.135 ;
        RECT  7.020 1.475 7.750 1.735 ;
        RECT  7.410 1.975 7.670 2.235 ;
        RECT  7.295 2.585 7.455 3.100 ;
        RECT  7.020 2.940 7.295 3.100 ;
        RECT  7.130 0.950 7.290 1.215 ;
        RECT  6.935 1.475 7.020 2.535 ;
        RECT  6.970 2.940 7.020 3.200 ;
        RECT  6.760 2.890 6.970 3.200 ;
        RECT  6.860 0.600 6.935 2.535 ;
        RECT  6.775 0.600 6.860 1.650 ;
        RECT  6.755 2.375 6.860 2.535 ;
        RECT  6.440 0.600 6.775 0.900 ;
        RECT  4.580 2.890 6.760 3.100 ;
        RECT  6.495 2.375 6.755 2.635 ;
        RECT  6.535 1.815 6.660 2.075 ;
        RECT  6.375 1.105 6.535 2.075 ;
        RECT  5.020 2.475 6.495 2.635 ;
        RECT  6.390 0.600 6.440 0.890 ;
        RECT  4.670 0.720 6.390 0.880 ;
        RECT  4.220 1.105 6.375 1.265 ;
        RECT  5.190 1.915 6.375 2.075 ;
        RECT  6.010 1.450 6.170 1.720 ;
        RECT  4.580 1.450 6.010 1.610 ;
        RECT  4.980 1.795 5.190 2.075 ;
        RECT  4.760 2.375 5.020 2.635 ;
        RECT  4.930 1.795 4.980 1.955 ;
        RECT  4.460 0.720 4.670 0.910 ;
        RECT  4.420 1.450 4.580 3.100 ;
        RECT  4.410 0.750 4.460 0.910 ;
        RECT  3.915 2.890 4.420 3.050 ;
        RECT  3.865 1.715 4.225 1.975 ;
        RECT  4.060 0.585 4.220 1.265 ;
        RECT  1.875 0.585 4.060 0.745 ;
        RECT  3.755 2.890 3.915 3.100 ;
        RECT  3.705 1.015 3.865 2.425 ;
        RECT  1.840 2.940 3.755 3.100 ;
        RECT  3.110 1.015 3.705 1.175 ;
        RECT  3.525 2.265 3.705 2.425 ;
        RECT  3.365 2.265 3.525 2.665 ;
        RECT  3.185 1.620 3.510 1.880 ;
        RECT  3.025 1.355 3.185 2.695 ;
        RECT  2.905 1.355 3.025 1.515 ;
        RECT  2.805 2.535 3.025 2.695 ;
        RECT  2.745 0.925 2.905 1.515 ;
        RECT  2.265 0.925 2.745 1.085 ;
        RECT  1.780 0.585 1.875 1.290 ;
        RECT  1.680 2.530 1.840 3.100 ;
        RECT  1.780 2.185 1.805 2.345 ;
        RECT  1.715 0.585 1.780 2.345 ;
        RECT  1.620 1.080 1.715 2.345 ;
        RECT  1.305 2.530 1.680 2.690 ;
        RECT  1.545 2.185 1.620 2.345 ;
        RECT  1.305 1.715 1.430 1.975 ;
        RECT  1.145 1.115 1.305 2.690 ;
        RECT  0.945 1.115 1.145 1.275 ;
        RECT  0.895 2.465 1.145 2.690 ;
        RECT  0.685 0.675 0.945 1.275 ;
        RECT  0.635 2.465 0.895 3.085 ;
    END
END TLATNTSCAX6

MACRO TLATNTSCAX4
    CLASS CORE ;
    FOREIGN TLATNTSCAX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.295 1.795 1.455 ;
        RECT  1.505 1.290 1.715 1.950 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.695 2.115 7.795 2.715 ;
        RECT  7.690 1.515 7.695 2.715 ;
        RECT  7.535 0.945 7.690 2.715 ;
        RECT  7.485 0.945 7.535 2.585 ;
        RECT  7.450 0.945 7.485 2.455 ;
        RECT  7.415 0.945 7.450 1.205 ;
        END
        ANTENNADIFFAREA     0.7410 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 1.700 2.235 2.140 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.765 0.370 2.045 ;
        RECT  0.125 1.575 0.345 2.145 ;
        END
        ANTENNAGATEAREA     0.2652 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.225 -0.250 8.740 0.250 ;
        RECT  7.965 -0.250 8.225 0.405 ;
        RECT  7.125 -0.250 7.965 0.250 ;
        RECT  6.865 -0.250 7.125 0.405 ;
        RECT  6.435 -0.250 6.865 0.250 ;
        RECT  6.175 -0.250 6.435 0.405 ;
        RECT  4.895 -0.250 6.175 0.250 ;
        RECT  4.635 -0.250 4.895 0.405 ;
        RECT  2.985 -0.250 4.635 0.250 ;
        RECT  2.385 -0.250 2.985 0.405 ;
        RECT  1.320 -0.250 2.385 0.250 ;
        RECT  0.720 -0.250 1.320 0.405 ;
        RECT  0.000 -0.250 0.720 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.615 3.440 8.740 3.940 ;
        RECT  8.355 2.275 8.615 3.940 ;
        RECT  6.840 3.440 8.355 3.940 ;
        RECT  6.580 2.945 6.840 3.940 ;
        RECT  5.245 3.440 6.580 3.940 ;
        RECT  4.985 3.285 5.245 3.940 ;
        RECT  3.525 3.440 4.985 3.940 ;
        RECT  3.265 3.285 3.525 3.940 ;
        RECT  1.440 3.440 3.265 3.940 ;
        RECT  1.180 2.955 1.440 3.940 ;
        RECT  0.385 3.440 1.180 3.940 ;
        RECT  0.125 2.800 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.315 1.740 8.575 2.000 ;
        RECT  8.160 1.840 8.315 2.000 ;
        RECT  8.000 1.840 8.160 3.215 ;
        RECT  7.880 0.605 8.040 1.640 ;
        RECT  7.265 3.055 8.000 3.215 ;
        RECT  5.770 0.605 7.880 0.765 ;
        RECT  7.105 1.375 7.265 3.215 ;
        RECT  6.290 2.585 7.105 2.745 ;
        RECT  6.765 1.055 6.925 2.185 ;
        RECT  6.125 1.055 6.765 1.215 ;
        RECT  6.505 2.025 6.765 2.185 ;
        RECT  5.770 1.475 6.585 1.735 ;
        RECT  6.245 1.955 6.505 2.215 ;
        RECT  6.130 2.585 6.290 3.100 ;
        RECT  5.805 2.940 6.130 3.100 ;
        RECT  5.965 0.950 6.125 1.215 ;
        RECT  5.545 2.940 5.805 3.200 ;
        RECT  5.610 0.605 5.770 2.635 ;
        RECT  5.225 0.605 5.610 0.920 ;
        RECT  5.605 2.475 5.610 2.635 ;
        RECT  5.345 2.475 5.605 2.735 ;
        RECT  4.835 2.940 5.545 3.100 ;
        RECT  5.025 1.235 5.420 1.495 ;
        RECT  4.385 2.475 5.345 2.635 ;
        RECT  3.775 0.760 5.225 0.920 ;
        RECT  4.865 1.105 5.025 1.905 ;
        RECT  3.595 1.105 4.865 1.265 ;
        RECT  4.555 1.745 4.865 1.905 ;
        RECT  3.915 2.850 4.835 3.100 ;
        RECT  4.295 1.745 4.555 2.005 ;
        RECT  4.125 2.375 4.385 2.635 ;
        RECT  3.915 1.450 4.050 1.610 ;
        RECT  3.755 1.450 3.915 3.100 ;
        RECT  1.840 2.855 3.755 3.015 ;
        RECT  3.435 0.585 3.595 1.265 ;
        RECT  3.255 1.705 3.545 1.965 ;
        RECT  1.325 0.585 3.435 0.745 ;
        RECT  3.095 0.985 3.255 2.425 ;
        RECT  2.500 0.985 3.095 1.145 ;
        RECT  2.925 2.265 3.095 2.425 ;
        RECT  2.765 2.265 2.925 2.665 ;
        RECT  2.580 1.620 2.910 1.880 ;
        RECT  2.420 1.330 2.580 2.635 ;
        RECT  2.150 1.330 2.420 1.490 ;
        RECT  2.205 2.375 2.420 2.635 ;
        RECT  1.990 0.925 2.150 1.490 ;
        RECT  1.715 0.925 1.990 1.085 ;
        RECT  1.680 2.565 1.840 3.015 ;
        RECT  0.895 2.565 1.680 2.725 ;
        RECT  1.165 0.585 1.325 2.115 ;
        RECT  1.155 1.955 1.165 2.115 ;
        RECT  0.995 1.955 1.155 2.255 ;
        RECT  0.875 1.485 0.985 1.750 ;
        RECT  0.795 2.565 0.895 3.060 ;
        RECT  0.725 1.070 0.875 1.750 ;
        RECT  0.725 2.450 0.795 3.060 ;
        RECT  0.715 1.070 0.725 3.060 ;
        RECT  0.385 1.070 0.715 1.230 ;
        RECT  0.635 1.485 0.715 3.060 ;
        RECT  0.565 1.485 0.635 2.610 ;
        RECT  0.125 0.630 0.385 1.230 ;
    END
END TLATNTSCAX4

MACRO TLATNTSCAX3
    CLASS CORE ;
    FOREIGN TLATNTSCAX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.295 1.795 1.455 ;
        RECT  1.505 1.290 1.715 1.950 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.345 2.275 6.395 2.875 ;
        RECT  6.345 0.975 6.375 1.235 ;
        RECT  6.135 0.975 6.345 2.875 ;
        RECT  6.115 0.975 6.135 2.585 ;
        RECT  6.105 1.355 6.115 2.585 ;
        END
        ANTENNADIFFAREA     0.6118 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 1.700 2.375 2.025 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.765 0.370 2.045 ;
        RECT  0.125 1.575 0.345 2.145 ;
        END
        ANTENNAGATEAREA     0.2158 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.925 -0.250 7.360 0.250 ;
        RECT  6.665 -0.250 6.925 0.405 ;
        RECT  5.815 -0.250 6.665 0.250 ;
        RECT  5.555 -0.250 5.815 0.405 ;
        RECT  5.005 -0.250 5.555 0.250 ;
        RECT  4.745 -0.250 5.005 0.405 ;
        RECT  2.925 -0.250 4.745 0.250 ;
        RECT  2.325 -0.250 2.925 0.405 ;
        RECT  1.275 -0.250 2.325 0.250 ;
        RECT  1.015 -0.250 1.275 0.405 ;
        RECT  0.000 -0.250 1.015 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.215 3.440 7.360 3.940 ;
        RECT  6.955 2.465 7.215 3.940 ;
        RECT  5.495 3.440 6.955 3.940 ;
        RECT  4.895 2.945 5.495 3.940 ;
        RECT  3.075 3.440 4.895 3.940 ;
        RECT  2.815 3.285 3.075 3.940 ;
        RECT  1.445 3.440 2.815 3.940 ;
        RECT  1.185 2.745 1.445 3.940 ;
        RECT  0.385 3.440 1.185 3.940 ;
        RECT  0.125 2.825 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.785 1.890 7.045 2.150 ;
        RECT  6.750 1.400 6.800 1.660 ;
        RECT  6.750 1.990 6.785 2.150 ;
        RECT  6.590 0.590 6.750 1.660 ;
        RECT  6.590 1.990 6.750 3.215 ;
        RECT  4.650 0.590 6.590 0.750 ;
        RECT  6.540 1.400 6.590 1.660 ;
        RECT  5.880 3.055 6.590 3.215 ;
        RECT  5.720 1.400 5.880 3.215 ;
        RECT  4.480 2.600 5.720 2.760 ;
        RECT  5.380 1.070 5.540 2.170 ;
        RECT  4.965 1.070 5.380 1.230 ;
        RECT  5.105 2.010 5.380 2.170 ;
        RECT  4.650 1.435 5.200 1.695 ;
        RECT  4.845 2.010 5.105 2.315 ;
        RECT  4.730 2.155 4.845 2.315 ;
        RECT  4.470 2.155 4.730 2.415 ;
        RECT  4.490 0.590 4.650 1.950 ;
        RECT  4.035 0.590 4.490 0.770 ;
        RECT  3.975 1.790 4.490 1.950 ;
        RECT  4.320 2.600 4.480 3.040 ;
        RECT  4.310 2.880 4.320 3.040 ;
        RECT  4.050 2.880 4.310 3.140 ;
        RECT  4.180 1.345 4.280 1.605 ;
        RECT  4.020 1.015 4.180 1.605 ;
        RECT  3.535 2.880 4.050 3.090 ;
        RECT  3.775 0.560 4.035 0.820 ;
        RECT  3.565 1.015 4.020 1.175 ;
        RECT  3.815 1.790 3.975 2.655 ;
        RECT  3.715 2.055 3.815 2.655 ;
        RECT  3.535 1.395 3.795 1.555 ;
        RECT  3.405 0.585 3.565 1.175 ;
        RECT  3.375 1.395 3.535 3.090 ;
        RECT  1.325 0.585 3.405 0.745 ;
        RECT  2.635 2.930 3.375 3.090 ;
        RECT  3.035 0.985 3.195 2.735 ;
        RECT  2.345 0.985 3.035 1.145 ;
        RECT  2.285 2.575 3.035 2.735 ;
        RECT  2.555 1.330 2.715 2.375 ;
        RECT  2.475 2.930 2.635 3.255 ;
        RECT  2.150 1.330 2.555 1.490 ;
        RECT  2.240 2.215 2.555 2.375 ;
        RECT  1.810 3.095 2.475 3.255 ;
        RECT  2.125 2.575 2.285 2.915 ;
        RECT  1.990 0.925 2.150 1.490 ;
        RECT  2.025 2.755 2.125 2.915 ;
        RECT  1.685 0.925 1.990 1.085 ;
        RECT  1.650 2.400 1.810 3.255 ;
        RECT  0.895 2.400 1.650 2.560 ;
        RECT  1.165 0.585 1.325 2.115 ;
        RECT  1.115 1.955 1.165 2.115 ;
        RECT  0.955 1.955 1.115 2.215 ;
        RECT  0.725 1.490 0.985 1.750 ;
        RECT  0.725 2.400 0.895 3.085 ;
        RECT  0.720 1.490 0.725 3.085 ;
        RECT  0.635 1.130 0.720 3.085 ;
        RECT  0.565 1.130 0.635 2.560 ;
        RECT  0.560 1.130 0.565 1.650 ;
        RECT  0.385 1.130 0.560 1.290 ;
        RECT  0.125 0.690 0.385 1.290 ;
    END
END TLATNTSCAX3

MACRO TLATNTSCAX2
    CLASS CORE ;
    FOREIGN TLATNTSCAX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.275 1.745 1.535 ;
        RECT  1.505 1.275 1.715 1.830 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.055 2.030 6.315 3.120 ;
        RECT  5.940 2.030 6.055 2.190 ;
        RECT  5.780 0.970 5.940 2.190 ;
        RECT  5.575 0.970 5.780 1.230 ;
        END
        ANTENNADIFFAREA     0.6062 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 1.825 2.380 2.035 ;
        RECT  2.175 1.755 2.230 2.035 ;
        RECT  1.965 1.700 2.175 2.035 ;
        RECT  1.940 1.825 1.965 2.035 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.765 0.370 2.045 ;
        RECT  0.125 1.575 0.345 2.145 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 -0.250 6.440 0.250 ;
        RECT  6.055 -0.250 6.315 0.405 ;
        RECT  5.295 -0.250 6.055 0.250 ;
        RECT  4.575 -0.250 5.295 0.405 ;
        RECT  2.925 -0.250 4.575 0.250 ;
        RECT  2.325 -0.250 2.925 0.405 ;
        RECT  1.275 -0.250 2.325 0.250 ;
        RECT  0.935 -0.250 1.275 0.405 ;
        RECT  0.675 -0.250 0.935 0.755 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.455 3.440 6.440 3.940 ;
        RECT  5.195 3.285 5.455 3.940 ;
        RECT  3.075 3.440 5.195 3.940 ;
        RECT  2.815 3.285 3.075 3.940 ;
        RECT  1.495 3.440 2.815 3.940 ;
        RECT  1.235 2.860 1.495 3.940 ;
        RECT  0.410 3.440 1.235 3.940 ;
        RECT  0.150 2.905 0.410 3.940 ;
        RECT  0.000 3.440 0.150 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.120 0.595 6.280 1.735 ;
        RECT  4.415 0.595 6.120 0.755 ;
        RECT  5.440 1.555 5.600 3.095 ;
        RECT  4.375 2.935 5.440 3.095 ;
        RECT  5.100 1.070 5.260 2.075 ;
        RECT  4.855 1.070 5.100 1.230 ;
        RECT  4.970 1.915 5.100 2.075 ;
        RECT  4.760 1.915 4.970 2.215 ;
        RECT  4.415 1.455 4.920 1.715 ;
        RECT  4.595 0.970 4.855 1.230 ;
        RECT  4.600 1.915 4.760 2.590 ;
        RECT  4.255 0.595 4.415 2.420 ;
        RECT  4.215 2.935 4.375 3.215 ;
        RECT  3.955 0.610 4.255 0.820 ;
        RECT  3.970 2.260 4.255 2.420 ;
        RECT  3.525 3.055 4.215 3.215 ;
        RECT  3.915 1.005 4.075 2.075 ;
        RECT  3.710 2.260 3.970 2.860 ;
        RECT  3.695 0.560 3.955 0.820 ;
        RECT  3.470 1.005 3.915 1.165 ;
        RECT  3.765 1.815 3.915 2.075 ;
        RECT  3.525 1.355 3.730 1.515 ;
        RECT  3.365 1.355 3.525 3.215 ;
        RECT  3.310 0.585 3.470 1.165 ;
        RECT  2.625 2.935 3.365 3.095 ;
        RECT  1.325 0.585 3.310 0.745 ;
        RECT  3.080 1.835 3.180 2.095 ;
        RECT  2.920 1.000 3.080 2.735 ;
        RECT  2.305 1.000 2.920 1.160 ;
        RECT  2.285 2.575 2.920 2.735 ;
        RECT  2.560 1.345 2.720 2.375 ;
        RECT  2.465 2.935 2.625 3.260 ;
        RECT  2.460 1.345 2.560 1.615 ;
        RECT  2.175 2.215 2.560 2.375 ;
        RECT  1.835 3.100 2.465 3.260 ;
        RECT  2.120 1.345 2.460 1.505 ;
        RECT  2.125 2.575 2.285 2.920 ;
        RECT  2.025 2.760 2.125 2.920 ;
        RECT  1.960 0.925 2.120 1.505 ;
        RECT  1.685 0.925 1.960 1.085 ;
        RECT  1.675 2.485 1.835 3.260 ;
        RECT  0.920 2.485 1.675 2.645 ;
        RECT  1.165 0.585 1.325 2.135 ;
        RECT  1.050 1.975 1.165 2.135 ;
        RECT  0.890 1.975 1.050 2.235 ;
        RECT  0.765 1.490 0.985 1.750 ;
        RECT  0.710 2.485 0.920 3.160 ;
        RECT  0.710 1.060 0.765 1.750 ;
        RECT  0.660 1.060 0.710 3.160 ;
        RECT  0.605 1.060 0.660 2.645 ;
        RECT  0.385 1.060 0.605 1.220 ;
        RECT  0.550 1.590 0.605 2.645 ;
        RECT  0.125 0.960 0.385 1.220 ;
    END
END TLATNTSCAX2

MACRO TLATNCAX20
    CLASS CORE ;
    FOREIGN TLATNCAX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.625 1.755 17.730 2.690 ;
        RECT  17.470 0.705 17.625 2.690 ;
        RECT  16.650 0.705 17.470 2.355 ;
        RECT  16.225 0.705 16.650 2.650 ;
        RECT  15.415 0.705 16.225 1.305 ;
        RECT  15.600 2.045 16.225 2.650 ;
        RECT  15.340 2.045 15.600 3.115 ;
        RECT  15.155 0.680 15.415 1.305 ;
        RECT  15.305 2.045 15.340 3.000 ;
        RECT  14.595 2.045 15.305 2.650 ;
        RECT  14.315 0.705 15.155 1.305 ;
        RECT  14.580 2.045 14.595 2.995 ;
        RECT  14.320 2.045 14.580 3.115 ;
        RECT  13.560 2.045 14.320 2.650 ;
        RECT  14.055 0.680 14.315 1.305 ;
        RECT  13.215 0.705 14.055 1.305 ;
        RECT  13.300 2.045 13.560 3.115 ;
        RECT  12.540 2.045 13.300 2.650 ;
        RECT  12.955 0.680 13.215 1.305 ;
        RECT  12.115 0.705 12.955 1.305 ;
        RECT  12.280 2.045 12.540 3.115 ;
        RECT  11.520 2.045 12.280 2.650 ;
        RECT  11.855 0.680 12.115 1.305 ;
        RECT  11.015 0.705 11.855 1.305 ;
        RECT  11.260 2.045 11.520 3.115 ;
        RECT  10.500 2.045 11.260 2.650 ;
        RECT  10.755 0.680 11.015 1.305 ;
        RECT  10.585 0.705 10.755 1.305 ;
        RECT  10.240 2.045 10.500 3.115 ;
        END
        ANTENNADIFFAREA     5.4785 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.415 1.810 1.675 ;
        RECT  1.550 1.415 1.765 2.090 ;
        RECT  1.505 1.515 1.550 1.990 ;
        END
        ANTENNAGATEAREA     0.3536 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.600 0.465 1.860 ;
        RECT  0.125 1.545 0.345 2.060 ;
        END
        ANTENNAGATEAREA     0.2691 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.970 -0.250 18.400 0.250 ;
        RECT  15.710 -0.250 15.970 0.405 ;
        RECT  14.865 -0.250 15.710 0.250 ;
        RECT  14.605 -0.250 14.865 0.405 ;
        RECT  13.765 -0.250 14.605 0.250 ;
        RECT  13.505 -0.250 13.765 0.405 ;
        RECT  12.665 -0.250 13.505 0.250 ;
        RECT  12.405 -0.250 12.665 0.405 ;
        RECT  11.565 -0.250 12.405 0.250 ;
        RECT  11.305 -0.250 11.565 0.405 ;
        RECT  10.445 -0.250 11.305 0.250 ;
        RECT  10.185 -0.250 10.445 0.405 ;
        RECT  9.435 -0.250 10.185 0.250 ;
        RECT  9.175 -0.250 9.435 0.405 ;
        RECT  8.400 -0.250 9.175 0.250 ;
        RECT  8.140 -0.250 8.400 0.405 ;
        RECT  7.355 -0.250 8.140 0.250 ;
        RECT  7.095 -0.250 7.355 0.405 ;
        RECT  6.260 -0.250 7.095 0.250 ;
        RECT  6.000 -0.250 6.260 0.405 ;
        RECT  5.195 -0.250 6.000 0.250 ;
        RECT  4.475 -0.250 5.195 0.405 ;
        RECT  3.450 -0.250 4.475 0.250 ;
        RECT  3.190 -0.250 3.450 0.405 ;
        RECT  1.730 -0.250 3.190 0.250 ;
        RECT  0.790 -0.250 1.730 0.405 ;
        RECT  0.000 -0.250 0.790 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.270 3.440 18.400 3.940 ;
        RECT  18.010 2.085 18.270 3.940 ;
        RECT  17.360 3.440 18.010 3.940 ;
        RECT  17.185 3.285 17.360 3.940 ;
        RECT  16.925 2.570 17.185 3.940 ;
        RECT  16.110 3.440 16.925 3.940 ;
        RECT  15.850 2.895 16.110 3.940 ;
        RECT  15.090 3.440 15.850 3.940 ;
        RECT  14.830 2.895 15.090 3.940 ;
        RECT  14.070 3.440 14.830 3.940 ;
        RECT  13.810 2.895 14.070 3.940 ;
        RECT  13.050 3.440 13.810 3.940 ;
        RECT  12.790 2.895 13.050 3.940 ;
        RECT  12.030 3.440 12.790 3.940 ;
        RECT  11.770 2.895 12.030 3.940 ;
        RECT  11.010 3.440 11.770 3.940 ;
        RECT  10.750 2.895 11.010 3.940 ;
        RECT  9.990 3.440 10.750 3.940 ;
        RECT  9.730 2.105 9.990 3.940 ;
        RECT  8.970 3.440 9.730 3.940 ;
        RECT  8.710 2.510 8.970 3.940 ;
        RECT  7.950 3.440 8.710 3.940 ;
        RECT  7.690 2.510 7.950 3.940 ;
        RECT  6.930 3.440 7.690 3.940 ;
        RECT  6.670 2.300 6.930 3.940 ;
        RECT  5.250 3.440 6.670 3.940 ;
        RECT  4.990 3.285 5.250 3.940 ;
        RECT  3.465 3.440 4.990 3.940 ;
        RECT  3.205 3.285 3.465 3.940 ;
        RECT  1.660 3.440 3.205 3.940 ;
        RECT  0.720 3.285 1.660 3.940 ;
        RECT  0.000 3.440 0.720 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.365 1.545 15.895 1.795 ;
        RECT  10.205 1.025 10.365 1.795 ;
        RECT  9.960 1.025 10.205 1.185 ;
        RECT  9.545 0.605 9.960 1.185 ;
        RECT  9.480 0.605 9.545 2.350 ;
        RECT  9.385 0.605 9.480 3.045 ;
        RECT  7.625 0.605 9.385 1.185 ;
        RECT  9.220 2.015 9.385 3.045 ;
        RECT  8.460 2.015 9.220 2.330 ;
        RECT  6.745 1.435 9.180 1.695 ;
        RECT  8.200 2.015 8.460 3.070 ;
        RECT  7.440 2.015 8.200 2.330 ;
        RECT  7.180 2.015 7.440 2.955 ;
        RECT  6.745 0.925 6.810 1.185 ;
        RECT  6.590 0.925 6.745 1.695 ;
        RECT  6.585 0.925 6.590 2.075 ;
        RECT  6.550 0.925 6.585 1.185 ;
        RECT  6.430 1.535 6.585 2.075 ;
        RECT  6.110 1.915 6.430 2.075 ;
        RECT  6.020 0.585 6.180 1.715 ;
        RECT  5.850 1.915 6.110 2.910 ;
        RECT  4.355 0.585 6.020 0.745 ;
        RECT  5.840 1.915 5.850 2.075 ;
        RECT  5.680 0.925 5.840 2.075 ;
        RECT  5.475 0.925 5.680 1.085 ;
        RECT  5.340 1.265 5.500 2.940 ;
        RECT  4.200 2.780 5.340 2.940 ;
        RECT  4.995 1.135 5.155 2.115 ;
        RECT  4.695 1.135 4.995 1.295 ;
        RECT  4.765 1.955 4.995 2.115 ;
        RECT  4.410 1.480 4.800 1.740 ;
        RECT  4.665 1.955 4.765 2.215 ;
        RECT  4.535 1.035 4.695 1.295 ;
        RECT  4.505 1.955 4.665 2.590 ;
        RECT  4.440 2.195 4.505 2.590 ;
        RECT  4.355 1.480 4.410 1.775 ;
        RECT  4.195 0.585 4.355 1.775 ;
        RECT  4.050 2.190 4.200 3.105 ;
        RECT  4.190 0.770 4.195 1.775 ;
        RECT  3.855 0.770 4.190 0.930 ;
        RECT  3.495 1.615 4.190 1.775 ;
        RECT  4.040 2.095 4.050 3.105 ;
        RECT  3.790 2.095 4.040 2.355 ;
        RECT  2.140 2.945 4.040 3.105 ;
        RECT  3.750 1.165 4.010 1.425 ;
        RECT  3.595 0.705 3.855 0.965 ;
        RECT  3.590 2.555 3.855 2.765 ;
        RECT  3.120 1.215 3.750 1.375 ;
        RECT  2.590 0.780 3.595 0.940 ;
        RECT  3.495 2.555 3.590 2.735 ;
        RECT  3.335 1.615 3.495 2.735 ;
        RECT  2.605 2.440 3.335 2.600 ;
        RECT  2.960 1.215 3.120 2.010 ;
        RECT  2.775 1.850 2.960 2.010 ;
        RECT  2.175 1.850 2.775 2.110 ;
        RECT  2.540 1.345 2.760 1.605 ;
        RECT  2.345 2.390 2.605 2.650 ;
        RECT  2.330 0.730 2.590 0.990 ;
        RECT  2.160 1.340 2.540 1.605 ;
        RECT  2.135 1.950 2.175 2.110 ;
        RECT  2.150 1.340 2.160 1.500 ;
        RECT  1.990 0.680 2.150 1.500 ;
        RECT  1.980 2.625 2.140 3.105 ;
        RECT  1.975 1.950 2.135 2.435 ;
        RECT  0.880 0.680 1.990 0.840 ;
        RECT  0.880 2.625 1.980 2.785 ;
        RECT  1.335 2.275 1.975 2.435 ;
        RECT  1.325 2.130 1.335 2.435 ;
        RECT  1.320 1.080 1.325 2.435 ;
        RECT  1.165 1.030 1.320 2.435 ;
        RECT  1.160 1.030 1.165 1.290 ;
        RECT  1.075 2.130 1.165 2.435 ;
        RECT  0.880 1.490 0.985 1.750 ;
        RECT  0.720 0.680 0.880 2.785 ;
        RECT  0.385 1.130 0.720 1.290 ;
        RECT  0.385 2.255 0.720 2.455 ;
        RECT  0.125 0.690 0.385 1.290 ;
        RECT  0.125 2.255 0.385 3.195 ;
    END
END TLATNCAX20

MACRO TLATNCAX16
    CLASS CORE ;
    FOREIGN TLATNCAX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.100 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.495 0.705 15.515 2.175 ;
        RECT  15.460 0.705 15.495 2.345 ;
        RECT  15.200 0.705 15.460 2.640 ;
        RECT  14.540 0.705 15.200 2.475 ;
        RECT  14.115 0.705 14.540 2.640 ;
        RECT  13.300 0.705 14.115 1.305 ;
        RECT  13.490 2.035 14.115 2.640 ;
        RECT  13.230 2.035 13.490 3.105 ;
        RECT  13.040 0.680 13.300 1.305 ;
        RECT  12.470 2.035 13.230 2.640 ;
        RECT  12.200 0.705 13.040 1.305 ;
        RECT  12.210 2.035 12.470 3.105 ;
        RECT  11.450 2.035 12.210 2.640 ;
        RECT  11.940 0.680 12.200 1.305 ;
        RECT  11.100 0.705 11.940 1.305 ;
        RECT  11.190 2.035 11.450 3.105 ;
        RECT  11.165 2.035 11.190 2.995 ;
        RECT  10.455 2.035 11.165 2.640 ;
        RECT  10.840 0.680 11.100 1.305 ;
        RECT  10.000 0.705 10.840 1.305 ;
        RECT  10.430 2.035 10.455 2.995 ;
        RECT  10.170 2.035 10.430 3.105 ;
        RECT  9.410 2.035 10.170 2.640 ;
        RECT  9.740 0.680 10.000 1.305 ;
        RECT  9.570 0.705 9.740 1.305 ;
        RECT  9.150 2.035 9.410 3.105 ;
        END
        ANTENNADIFFAREA     4.8346 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.415 1.815 1.675 ;
        RECT  1.555 1.415 1.770 2.090 ;
        RECT  1.505 1.700 1.555 1.990 ;
        END
        ANTENNAGATEAREA     0.2574 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.600 0.465 1.860 ;
        RECT  0.125 1.545 0.345 2.060 ;
        END
        ANTENNAGATEAREA     0.2158 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.850 -0.250 16.100 0.250 ;
        RECT  13.590 -0.250 13.850 0.405 ;
        RECT  12.750 -0.250 13.590 0.250 ;
        RECT  12.490 -0.250 12.750 0.405 ;
        RECT  11.650 -0.250 12.490 0.250 ;
        RECT  11.390 -0.250 11.650 0.405 ;
        RECT  10.550 -0.250 11.390 0.250 ;
        RECT  10.290 -0.250 10.550 0.405 ;
        RECT  9.450 -0.250 10.290 0.250 ;
        RECT  9.190 -0.250 9.450 0.405 ;
        RECT  8.350 -0.250 9.190 0.250 ;
        RECT  8.090 -0.250 8.350 0.405 ;
        RECT  7.245 -0.250 8.090 0.250 ;
        RECT  6.985 -0.250 7.245 0.405 ;
        RECT  6.190 -0.250 6.985 0.250 ;
        RECT  5.930 -0.250 6.190 0.405 ;
        RECT  5.085 -0.250 5.930 0.250 ;
        RECT  4.825 -0.250 5.085 0.405 ;
        RECT  3.995 -0.250 4.825 0.250 ;
        RECT  3.275 -0.250 3.995 0.405 ;
        RECT  1.730 -0.250 3.275 0.250 ;
        RECT  0.790 -0.250 1.730 0.405 ;
        RECT  0.000 -0.250 0.790 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.970 3.440 16.100 3.940 ;
        RECT  15.710 2.075 15.970 3.940 ;
        RECT  14.990 3.440 15.710 3.940 ;
        RECT  14.730 3.285 14.990 3.940 ;
        RECT  14.000 3.440 14.730 3.940 ;
        RECT  13.740 2.885 14.000 3.940 ;
        RECT  12.980 3.440 13.740 3.940 ;
        RECT  12.720 2.885 12.980 3.940 ;
        RECT  11.960 3.440 12.720 3.940 ;
        RECT  11.700 2.885 11.960 3.940 ;
        RECT  10.940 3.440 11.700 3.940 ;
        RECT  10.680 2.885 10.940 3.940 ;
        RECT  9.920 3.440 10.680 3.940 ;
        RECT  9.660 2.885 9.920 3.940 ;
        RECT  8.900 3.440 9.660 3.940 ;
        RECT  8.640 2.095 8.900 3.940 ;
        RECT  7.880 3.440 8.640 3.940 ;
        RECT  7.620 2.500 7.880 3.940 ;
        RECT  6.860 3.440 7.620 3.940 ;
        RECT  6.600 2.500 6.860 3.940 ;
        RECT  5.835 3.440 6.600 3.940 ;
        RECT  5.575 2.105 5.835 3.940 ;
        RECT  4.155 3.440 5.575 3.940 ;
        RECT  3.895 3.285 4.155 3.940 ;
        RECT  1.715 3.440 3.895 3.940 ;
        RECT  1.115 3.285 1.715 3.940 ;
        RECT  0.000 3.440 1.115 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.295 1.555 13.325 1.715 ;
        RECT  9.135 1.025 9.295 1.715 ;
        RECT  8.900 1.025 9.135 1.185 ;
        RECT  8.640 0.925 8.900 1.185 ;
        RECT  8.455 0.975 8.640 1.185 ;
        RECT  8.390 0.975 8.455 2.340 ;
        RECT  8.295 0.975 8.390 3.035 ;
        RECT  7.800 0.975 8.295 1.135 ;
        RECT  8.130 2.095 8.295 3.035 ;
        RECT  7.370 2.095 8.130 2.255 ;
        RECT  6.460 1.435 8.080 1.695 ;
        RECT  7.540 0.925 7.800 1.185 ;
        RECT  6.700 0.975 7.540 1.135 ;
        RECT  7.110 2.095 7.370 3.060 ;
        RECT  6.350 2.095 7.110 2.255 ;
        RECT  6.440 0.925 6.700 1.185 ;
        RECT  5.570 1.480 6.460 1.640 ;
        RECT  6.090 2.055 6.350 2.995 ;
        RECT  5.570 0.985 5.635 1.245 ;
        RECT  5.410 0.985 5.570 1.640 ;
        RECT  5.375 0.985 5.410 1.245 ;
        RECT  5.355 1.480 5.410 1.640 ;
        RECT  5.195 1.480 5.355 2.095 ;
        RECT  5.015 1.935 5.195 2.095 ;
        RECT  4.755 1.935 5.015 2.705 ;
        RECT  4.820 0.630 4.980 1.630 ;
        RECT  3.165 0.630 4.820 0.790 ;
        RECT  4.640 1.935 4.755 2.095 ;
        RECT  4.480 0.970 4.640 2.095 ;
        RECT  4.275 0.970 4.480 1.230 ;
        RECT  4.140 1.555 4.300 3.095 ;
        RECT  3.010 2.935 4.140 3.095 ;
        RECT  3.800 1.095 3.960 2.075 ;
        RECT  3.505 1.095 3.800 1.255 ;
        RECT  3.670 1.915 3.800 2.075 ;
        RECT  3.510 1.915 3.670 2.215 ;
        RECT  3.165 1.455 3.620 1.715 ;
        RECT  3.350 1.915 3.510 2.590 ;
        RECT  3.345 0.995 3.505 1.255 ;
        RECT  3.005 0.630 3.165 2.640 ;
        RECT  2.850 2.935 3.010 3.215 ;
        RECT  2.940 0.630 3.005 1.665 ;
        RECT  2.605 2.480 3.005 2.640 ;
        RECT  2.590 0.630 2.940 0.790 ;
        RECT  2.150 3.055 2.850 3.215 ;
        RECT  2.760 1.820 2.820 2.080 ;
        RECT  2.600 1.030 2.760 2.080 ;
        RECT  2.345 2.260 2.605 2.860 ;
        RECT  1.325 1.030 2.600 1.190 ;
        RECT  2.330 0.585 2.590 0.845 ;
        RECT  2.320 1.395 2.420 1.555 ;
        RECT  2.160 1.395 2.320 2.040 ;
        RECT  2.150 1.880 2.160 2.040 ;
        RECT  1.990 1.880 2.150 3.215 ;
        RECT  1.915 2.915 1.990 3.215 ;
        RECT  0.385 2.915 1.915 3.075 ;
        RECT  1.325 2.175 1.355 2.435 ;
        RECT  1.165 1.030 1.325 2.435 ;
        RECT  1.160 1.030 1.165 1.290 ;
        RECT  1.095 2.175 1.165 2.435 ;
        RECT  0.830 1.690 0.985 1.970 ;
        RECT  0.670 1.130 0.830 2.460 ;
        RECT  0.385 1.130 0.670 1.290 ;
        RECT  0.385 2.300 0.670 2.460 ;
        RECT  0.125 0.690 0.385 1.290 ;
        RECT  0.225 2.300 0.385 3.075 ;
        RECT  0.125 2.300 0.225 2.900 ;
    END
END TLATNCAX16

MACRO TLATNCAX12
    CLASS CORE ;
    FOREIGN TLATNCAX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.620 2.335 12.755 2.585 ;
        RECT  12.415 0.705 12.750 1.305 ;
        RECT  12.415 1.925 12.620 3.115 ;
        RECT  12.270 0.705 12.415 3.115 ;
        RECT  11.585 0.705 12.270 2.650 ;
        RECT  7.160 0.705 11.585 1.305 ;
        RECT  11.575 2.045 11.585 2.650 ;
        RECT  11.315 2.045 11.575 3.115 ;
        RECT  10.555 2.045 11.315 2.650 ;
        RECT  10.295 2.045 10.555 3.115 ;
        RECT  10.245 2.045 10.295 2.995 ;
        RECT  9.535 2.045 10.245 2.650 ;
        RECT  9.275 2.045 9.535 3.115 ;
        RECT  8.515 2.045 9.275 2.650 ;
        RECT  8.255 2.045 8.515 3.115 ;
        RECT  7.495 2.045 8.255 2.650 ;
        RECT  7.235 2.045 7.495 3.115 ;
        END
        ANTENNADIFFAREA     3.9040 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.415 1.810 1.675 ;
        RECT  1.550 1.415 1.765 2.090 ;
        RECT  1.505 1.700 1.550 1.990 ;
        END
        ANTENNAGATEAREA     0.2106 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.600 0.460 1.860 ;
        RECT  0.125 1.545 0.345 2.060 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.245 -0.250 12.880 0.250 ;
        RECT  11.985 -0.250 12.245 0.405 ;
        RECT  11.215 -0.250 11.985 0.250 ;
        RECT  10.955 -0.250 11.215 0.405 ;
        RECT  10.200 -0.250 10.955 0.250 ;
        RECT  9.940 -0.250 10.200 0.405 ;
        RECT  9.145 -0.250 9.940 0.250 ;
        RECT  8.885 -0.250 9.145 0.405 ;
        RECT  8.110 -0.250 8.885 0.250 ;
        RECT  7.850 -0.250 8.110 0.405 ;
        RECT  7.075 -0.250 7.850 0.250 ;
        RECT  6.815 -0.250 7.075 0.405 ;
        RECT  6.060 -0.250 6.815 0.250 ;
        RECT  5.800 -0.250 6.060 0.405 ;
        RECT  5.015 -0.250 5.800 0.250 ;
        RECT  4.755 -0.250 5.015 0.405 ;
        RECT  3.925 -0.250 4.755 0.250 ;
        RECT  3.205 -0.250 3.925 0.405 ;
        RECT  1.725 -0.250 3.205 0.250 ;
        RECT  0.785 -0.250 1.725 0.405 ;
        RECT  0.000 -0.250 0.785 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.085 3.440 12.880 3.940 ;
        RECT  11.825 2.895 12.085 3.940 ;
        RECT  11.065 3.440 11.825 3.940 ;
        RECT  10.805 2.895 11.065 3.940 ;
        RECT  10.045 3.440 10.805 3.940 ;
        RECT  9.785 2.895 10.045 3.940 ;
        RECT  9.025 3.440 9.785 3.940 ;
        RECT  8.765 2.895 9.025 3.940 ;
        RECT  8.005 3.440 8.765 3.940 ;
        RECT  7.745 2.895 8.005 3.940 ;
        RECT  6.985 3.440 7.745 3.940 ;
        RECT  6.725 2.105 6.985 3.940 ;
        RECT  5.965 3.440 6.725 3.940 ;
        RECT  5.705 2.575 5.965 3.940 ;
        RECT  4.085 3.440 5.705 3.940 ;
        RECT  3.825 3.285 4.085 3.940 ;
        RECT  1.710 3.440 3.825 3.940 ;
        RECT  1.110 3.285 1.710 3.940 ;
        RECT  0.000 3.440 1.110 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.565 1.555 11.085 1.715 ;
        RECT  6.540 0.925 6.565 1.715 ;
        RECT  6.475 0.925 6.540 2.350 ;
        RECT  6.380 0.925 6.475 3.045 ;
        RECT  6.305 0.925 6.380 1.185 ;
        RECT  6.215 2.105 6.380 3.045 ;
        RECT  5.525 1.025 6.305 1.185 ;
        RECT  5.455 2.195 6.215 2.355 ;
        RECT  5.915 1.440 6.135 1.700 ;
        RECT  5.590 1.435 5.915 1.700 ;
        RECT  5.430 1.435 5.590 1.945 ;
        RECT  5.265 0.925 5.525 1.185 ;
        RECT  5.195 2.195 5.455 3.135 ;
        RECT  4.945 1.785 5.430 1.945 ;
        RECT  4.960 1.420 5.010 1.580 ;
        RECT  4.800 0.595 4.960 1.580 ;
        RECT  4.685 1.785 4.945 3.045 ;
        RECT  3.095 0.595 4.800 0.755 ;
        RECT  4.750 1.420 4.800 1.580 ;
        RECT  4.570 1.785 4.685 1.945 ;
        RECT  4.410 0.970 4.570 1.945 ;
        RECT  4.205 0.970 4.410 1.230 ;
        RECT  4.070 1.555 4.230 3.095 ;
        RECT  3.005 2.935 4.070 3.095 ;
        RECT  3.730 1.095 3.890 2.075 ;
        RECT  3.435 1.095 3.730 1.255 ;
        RECT  3.600 1.915 3.730 2.075 ;
        RECT  3.440 1.915 3.600 2.215 ;
        RECT  3.095 1.455 3.550 1.715 ;
        RECT  3.280 1.915 3.440 2.590 ;
        RECT  3.275 0.995 3.435 1.255 ;
        RECT  2.935 0.595 3.095 2.640 ;
        RECT  2.845 2.935 3.005 3.215 ;
        RECT  2.325 0.650 2.935 0.810 ;
        RECT  2.600 2.480 2.935 2.640 ;
        RECT  2.145 3.055 2.845 3.215 ;
        RECT  2.595 1.030 2.755 2.080 ;
        RECT  2.340 2.260 2.600 2.860 ;
        RECT  1.325 1.030 2.595 1.190 ;
        RECT  2.575 1.820 2.595 2.080 ;
        RECT  2.365 1.375 2.415 1.535 ;
        RECT  2.335 1.375 2.365 1.540 ;
        RECT  2.175 1.375 2.335 2.040 ;
        RECT  2.155 1.375 2.175 1.535 ;
        RECT  2.145 1.880 2.175 2.040 ;
        RECT  1.985 1.880 2.145 3.215 ;
        RECT  1.910 2.915 1.985 3.215 ;
        RECT  0.385 2.915 1.910 3.075 ;
        RECT  1.325 2.240 1.355 2.500 ;
        RECT  1.165 1.030 1.325 2.500 ;
        RECT  1.155 1.030 1.165 1.295 ;
        RECT  1.095 2.240 1.165 2.500 ;
        RECT  0.830 1.690 0.985 1.970 ;
        RECT  0.670 1.060 0.830 2.460 ;
        RECT  0.385 1.060 0.670 1.220 ;
        RECT  0.385 2.300 0.670 2.460 ;
        RECT  0.125 0.960 0.385 1.220 ;
        RECT  0.225 2.300 0.385 3.075 ;
        RECT  0.125 2.300 0.225 2.900 ;
    END
END TLATNCAX12

MACRO TLATNCAX8
    CLASS CORE ;
    FOREIGN TLATNCAX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.800 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.675 0.665 13.680 2.405 ;
        RECT  13.650 0.665 13.675 3.000 ;
        RECT  13.390 0.665 13.650 3.195 ;
        RECT  13.280 0.665 13.390 2.810 ;
        RECT  8.350 0.665 13.280 1.065 ;
        RECT  13.005 2.005 13.280 2.810 ;
        RECT  12.080 2.005 13.005 2.405 ;
        RECT  11.680 2.005 12.080 3.195 ;
        RECT  11.625 2.005 11.680 2.995 ;
        RECT  10.455 2.005 11.625 2.405 ;
        RECT  10.440 2.005 10.455 2.995 ;
        RECT  10.040 2.005 10.440 3.195 ;
        RECT  8.870 2.005 10.040 2.405 ;
        RECT  8.470 2.005 8.870 3.045 ;
        RECT  8.405 2.335 8.470 2.585 ;
        END
        ANTENNADIFFAREA     2.5866 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.080 1.685 6.240 2.295 ;
        RECT  4.650 2.135 6.080 2.295 ;
        RECT  4.390 1.685 4.650 2.295 ;
        RECT  3.095 2.135 4.390 2.295 ;
        RECT  2.900 2.110 3.095 2.400 ;
        RECT  2.885 1.685 2.900 2.400 ;
        RECT  2.740 1.685 2.885 2.295 ;
        END
        ANTENNAGATEAREA     1.0140 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.565 1.065 1.825 ;
        RECT  0.585 1.565 0.795 1.990 ;
        RECT  0.465 1.565 0.585 1.825 ;
        END
        ANTENNAGATEAREA     0.8372 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.540 -0.250 13.800 0.250 ;
        RECT  13.280 -0.250 13.540 0.405 ;
        RECT  12.460 -0.250 13.280 0.250 ;
        RECT  12.200 -0.250 12.460 0.405 ;
        RECT  11.380 -0.250 12.200 0.250 ;
        RECT  11.120 -0.250 11.380 0.405 ;
        RECT  10.300 -0.250 11.120 0.250 ;
        RECT  10.040 -0.250 10.300 0.405 ;
        RECT  9.220 -0.250 10.040 0.250 ;
        RECT  8.960 -0.250 9.220 0.405 ;
        RECT  8.130 -0.250 8.960 0.250 ;
        RECT  7.870 -0.250 8.130 1.085 ;
        RECT  7.630 -0.250 7.870 0.285 ;
        RECT  7.280 -0.250 7.630 0.460 ;
        RECT  6.290 -0.250 7.280 0.250 ;
        RECT  6.030 -0.250 6.290 0.405 ;
        RECT  4.590 -0.250 6.030 0.250 ;
        RECT  4.330 -0.250 4.590 0.405 ;
        RECT  2.890 -0.250 4.330 0.250 ;
        RECT  2.630 -0.250 2.890 0.405 ;
        RECT  1.945 -0.250 2.630 0.250 ;
        RECT  1.685 -0.250 1.945 0.405 ;
        RECT  0.895 -0.250 1.685 0.250 ;
        RECT  0.635 -0.250 0.895 1.225 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.830 3.440 13.800 3.940 ;
        RECT  12.780 2.895 12.830 3.940 ;
        RECT  12.620 2.595 12.780 3.940 ;
        RECT  12.570 2.895 12.620 3.940 ;
        RECT  11.190 3.440 12.570 3.940 ;
        RECT  10.930 2.595 11.190 3.940 ;
        RECT  9.550 3.440 10.930 3.940 ;
        RECT  9.290 2.595 9.550 3.940 ;
        RECT  7.850 3.440 9.290 3.940 ;
        RECT  7.250 3.285 7.850 3.940 ;
        RECT  6.150 3.440 7.250 3.940 ;
        RECT  5.890 3.285 6.150 3.940 ;
        RECT  4.450 3.440 5.890 3.940 ;
        RECT  4.190 3.285 4.450 3.940 ;
        RECT  2.750 3.440 4.190 3.940 ;
        RECT  2.490 3.285 2.750 3.940 ;
        RECT  1.945 3.440 2.490 3.940 ;
        RECT  1.685 3.285 1.945 3.940 ;
        RECT  0.895 3.440 1.685 3.940 ;
        RECT  0.635 2.595 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.880 1.265 13.090 1.525 ;
        RECT  8.510 1.285 12.880 1.445 ;
        RECT  8.285 1.625 12.660 1.785 ;
        RECT  8.250 1.265 8.510 1.445 ;
        RECT  8.125 1.625 8.285 1.855 ;
        RECT  7.920 1.285 8.250 1.445 ;
        RECT  8.030 1.695 8.125 1.855 ;
        RECT  7.870 1.695 8.030 3.105 ;
        RECT  7.760 1.285 7.920 1.515 ;
        RECT  6.720 2.945 7.870 3.105 ;
        RECT  7.690 1.355 7.760 1.515 ;
        RECT  7.530 1.355 7.690 2.765 ;
        RECT  7.190 0.995 7.540 1.155 ;
        RECT  7.370 1.695 7.530 1.955 ;
        RECT  6.605 2.605 7.530 2.765 ;
        RECT  7.190 2.135 7.350 2.395 ;
        RECT  7.030 0.995 7.190 2.395 ;
        RECT  6.820 1.885 7.030 2.145 ;
        RECT  6.690 0.665 6.850 1.695 ;
        RECT  6.460 2.945 6.720 3.230 ;
        RECT  6.400 0.665 6.690 0.915 ;
        RECT  6.605 1.535 6.690 1.695 ;
        RECT  6.445 1.535 6.605 2.765 ;
        RECT  6.295 1.095 6.505 1.355 ;
        RECT  1.405 2.945 6.460 3.105 ;
        RECT  5.300 2.605 6.445 2.765 ;
        RECT  5.440 0.665 6.400 0.825 ;
        RECT  5.900 1.195 6.295 1.355 ;
        RECT  5.740 1.195 5.900 1.955 ;
        RECT  5.130 1.795 5.740 1.955 ;
        RECT  5.400 1.005 5.560 1.615 ;
        RECT  5.180 0.565 5.440 0.825 ;
        RECT  3.860 1.005 5.400 1.165 ;
        RECT  5.040 2.505 5.300 2.765 ;
        RECT  3.740 0.665 5.180 0.825 ;
        RECT  5.030 1.685 5.130 1.955 ;
        RECT  3.600 2.605 5.040 2.765 ;
        RECT  4.870 1.345 5.030 1.955 ;
        RECT  4.205 1.345 4.870 1.505 ;
        RECT  4.045 1.345 4.205 1.955 ;
        RECT  3.455 1.795 4.045 1.955 ;
        RECT  3.700 1.005 3.860 1.615 ;
        RECT  3.480 0.565 3.740 0.825 ;
        RECT  3.205 1.005 3.700 1.165 ;
        RECT  3.340 2.505 3.600 2.765 ;
        RECT  3.295 1.735 3.455 1.955 ;
        RECT  3.135 1.345 3.295 1.895 ;
        RECT  3.045 0.585 3.205 1.165 ;
        RECT  2.515 1.345 3.135 1.505 ;
        RECT  1.405 0.585 3.045 0.745 ;
        RECT  2.355 1.075 2.515 2.650 ;
        RECT  2.345 1.075 2.355 1.235 ;
        RECT  2.345 2.490 2.355 2.650 ;
        RECT  2.085 0.975 2.345 1.235 ;
        RECT  2.085 2.490 2.345 2.750 ;
        RECT  1.915 1.495 2.175 2.135 ;
        RECT  1.405 1.495 1.915 1.655 ;
        RECT  1.245 0.585 1.405 3.105 ;
        RECT  1.145 0.585 1.245 1.260 ;
        RECT  1.145 2.070 1.245 3.105 ;
        RECT  0.385 2.245 1.145 2.405 ;
        RECT  0.285 0.660 0.385 1.260 ;
        RECT  0.285 2.070 0.385 3.010 ;
        RECT  0.125 0.660 0.285 3.010 ;
    END
END TLATNCAX8

MACRO TLATNCAX6
    CLASS CORE ;
    FOREIGN TLATNCAX6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.155 0.695 8.160 2.585 ;
        RECT  7.895 0.695 8.155 3.105 ;
        RECT  7.860 0.695 7.895 2.435 ;
        RECT  6.225 0.695 7.860 0.995 ;
        RECT  7.485 1.700 7.860 2.435 ;
        RECT  6.535 2.135 7.485 2.435 ;
        RECT  6.235 2.135 6.535 3.105 ;
        RECT  6.105 2.335 6.235 2.585 ;
        END
        ANTENNADIFFAREA     1.4384 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.925 1.785 4.085 2.400 ;
        RECT  3.805 2.110 3.925 2.400 ;
        RECT  2.355 2.175 3.805 2.335 ;
        RECT  2.195 1.585 2.355 2.335 ;
        END
        ANTENNAGATEAREA     0.5044 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.515 0.865 1.990 ;
        END
        ANTENNAGATEAREA     0.4251 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.105 -0.250 8.280 0.250 ;
        RECT  7.845 -0.250 8.105 0.405 ;
        RECT  7.025 -0.250 7.845 0.250 ;
        RECT  6.765 -0.250 7.025 0.405 ;
        RECT  5.925 -0.250 6.765 0.250 ;
        RECT  5.765 -0.250 5.925 0.925 ;
        RECT  4.045 -0.250 5.765 0.250 ;
        RECT  3.785 -0.250 4.045 0.405 ;
        RECT  2.345 -0.250 3.785 0.250 ;
        RECT  1.175 -0.250 2.345 0.405 ;
        RECT  0.385 -0.250 1.175 0.250 ;
        RECT  0.125 -0.250 0.385 1.290 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.335 3.440 8.280 3.940 ;
        RECT  7.075 2.645 7.335 3.940 ;
        RECT  5.605 3.440 7.075 3.940 ;
        RECT  5.005 3.285 5.605 3.940 ;
        RECT  3.905 3.440 5.005 3.940 ;
        RECT  3.645 3.285 3.905 3.940 ;
        RECT  2.190 3.440 3.645 3.940 ;
        RECT  1.250 2.945 2.190 3.940 ;
        RECT  0.385 3.440 1.250 3.940 ;
        RECT  0.125 2.255 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.495 1.235 7.655 1.510 ;
        RECT  6.315 1.235 7.495 1.395 ;
        RECT  6.905 1.575 7.165 1.865 ;
        RECT  5.755 1.705 6.905 1.865 ;
        RECT  6.265 1.235 6.315 1.525 ;
        RECT  6.055 1.175 6.265 1.525 ;
        RECT  5.585 1.175 6.055 1.335 ;
        RECT  5.655 1.520 5.755 1.865 ;
        RECT  5.495 1.520 5.655 3.080 ;
        RECT  5.425 0.525 5.585 1.335 ;
        RECT  4.540 2.920 5.495 3.080 ;
        RECT  4.905 0.525 5.425 0.685 ;
        RECT  5.085 0.865 5.245 2.470 ;
        RECT  4.960 2.210 5.085 2.470 ;
        RECT  4.800 2.210 4.960 2.370 ;
        RECT  4.745 0.525 4.905 1.820 ;
        RECT  4.640 2.010 4.800 2.370 ;
        RECT  4.575 0.525 4.745 0.775 ;
        RECT  4.425 1.660 4.745 1.820 ;
        RECT  3.650 0.615 4.575 0.775 ;
        RECT  4.280 2.920 4.540 3.230 ;
        RECT  4.375 0.995 4.535 1.465 ;
        RECT  4.265 1.660 4.425 2.740 ;
        RECT  3.705 1.305 4.375 1.465 ;
        RECT  2.540 2.920 4.280 3.080 ;
        RECT  2.795 2.580 4.265 2.740 ;
        RECT  3.545 1.305 3.705 1.945 ;
        RECT  3.490 0.565 3.650 0.775 ;
        RECT  2.885 1.785 3.545 1.945 ;
        RECT  2.935 0.565 3.490 0.725 ;
        RECT  3.265 1.345 3.365 1.605 ;
        RECT  3.105 0.905 3.265 1.605 ;
        RECT  2.670 0.905 3.105 1.065 ;
        RECT  2.785 1.685 2.885 1.945 ;
        RECT  2.625 1.245 2.785 1.945 ;
        RECT  2.510 0.625 2.670 1.065 ;
        RECT  2.015 1.245 2.625 1.405 ;
        RECT  2.380 2.535 2.540 3.080 ;
        RECT  0.895 0.625 2.510 0.785 ;
        RECT  1.305 2.535 2.380 2.695 ;
        RECT  1.855 0.965 2.015 2.210 ;
        RECT  1.545 0.965 1.855 1.125 ;
        RECT  1.755 2.050 1.855 2.210 ;
        RECT  1.495 2.050 1.755 2.310 ;
        RECT  1.305 1.575 1.675 1.835 ;
        RECT  1.145 1.130 1.305 2.695 ;
        RECT  0.895 1.130 1.145 1.290 ;
        RECT  0.925 2.535 1.145 2.695 ;
        RECT  0.665 2.255 0.925 3.195 ;
        RECT  0.635 0.625 0.895 1.290 ;
    END
END TLATNCAX6

MACRO TLATNCAX4
    CLASS CORE ;
    FOREIGN TLATNCAX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.175 0.610 6.235 1.210 ;
        RECT  5.975 0.610 6.175 2.075 ;
        RECT  5.905 1.875 5.975 2.075 ;
        RECT  5.745 1.875 5.905 2.890 ;
        RECT  5.705 1.875 5.745 2.810 ;
        RECT  5.645 2.110 5.705 2.810 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.290 3.095 1.765 ;
        RECT  1.920 1.585 2.885 1.745 ;
        END
        ANTENNAGATEAREA     0.3796 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.570 0.415 2.000 ;
        END
        ANTENNAGATEAREA     0.2704 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 -0.250 6.900 0.250 ;
        RECT  6.515 -0.250 6.775 1.135 ;
        RECT  5.645 -0.250 6.515 0.250 ;
        RECT  5.485 -0.250 5.645 1.065 ;
        RECT  3.455 -0.250 5.485 0.250 ;
        RECT  3.195 -0.250 3.455 0.405 ;
        RECT  1.745 -0.250 3.195 0.250 ;
        RECT  1.485 -0.250 1.745 0.405 ;
        RECT  0.385 -0.250 1.485 0.250 ;
        RECT  0.125 -0.250 0.385 1.135 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.595 6.775 3.940 ;
        RECT  5.090 3.440 6.515 3.940 ;
        RECT  4.490 2.895 5.090 3.940 ;
        RECT  3.340 3.440 4.490 3.940 ;
        RECT  3.080 3.285 3.340 3.940 ;
        RECT  1.550 3.440 3.080 3.940 ;
        RECT  1.290 2.895 1.550 3.940 ;
        RECT  0.385 3.440 1.290 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.515 1.585 6.615 1.845 ;
        RECT  6.355 1.585 6.515 2.415 ;
        RECT  6.295 2.255 6.355 2.415 ;
        RECT  6.135 2.255 6.295 3.230 ;
        RECT  5.465 3.070 6.135 3.230 ;
        RECT  5.685 1.435 5.785 1.695 ;
        RECT  5.525 1.245 5.685 1.695 ;
        RECT  5.305 1.245 5.525 1.405 ;
        RECT  5.305 2.525 5.465 3.230 ;
        RECT  5.145 0.685 5.305 1.405 ;
        RECT  5.255 2.525 5.305 2.685 ;
        RECT  5.095 1.585 5.255 2.685 ;
        RECT  4.575 0.685 5.145 0.845 ;
        RECT  4.115 2.525 5.095 2.685 ;
        RECT  4.915 1.025 4.965 1.285 ;
        RECT  4.755 1.025 4.915 2.115 ;
        RECT  4.590 1.955 4.755 2.115 ;
        RECT  4.330 1.955 4.590 2.215 ;
        RECT  4.415 0.685 4.575 1.775 ;
        RECT  4.035 0.795 4.415 1.055 ;
        RECT  3.775 1.615 4.415 1.775 ;
        RECT  3.960 1.955 4.330 2.115 ;
        RECT  3.435 1.235 4.145 1.395 ;
        RECT  3.955 2.525 4.115 3.075 ;
        RECT  2.605 0.845 4.035 1.005 ;
        RECT  3.910 2.915 3.955 3.075 ;
        RECT  3.650 2.915 3.910 3.105 ;
        RECT  3.615 1.615 3.775 2.735 ;
        RECT  1.985 2.915 3.650 3.075 ;
        RECT  2.490 2.575 3.615 2.735 ;
        RECT  3.275 1.235 3.435 2.135 ;
        RECT  2.660 1.975 3.275 2.135 ;
        RECT  2.135 1.245 2.660 1.405 ;
        RECT  2.400 1.975 2.660 2.235 ;
        RECT  2.345 0.720 2.605 1.005 ;
        RECT  2.230 2.475 2.490 2.735 ;
        RECT  1.740 2.035 2.400 2.195 ;
        RECT  1.975 0.695 2.135 1.405 ;
        RECT  1.825 2.540 1.985 3.075 ;
        RECT  0.925 0.695 1.975 0.855 ;
        RECT  0.925 2.540 1.825 2.700 ;
        RECT  1.580 1.135 1.740 2.195 ;
        RECT  1.325 1.135 1.580 1.295 ;
        RECT  1.210 2.035 1.580 2.195 ;
        RECT  0.825 1.585 1.400 1.845 ;
        RECT  1.065 1.035 1.325 1.295 ;
        RECT  0.950 2.035 1.210 2.295 ;
        RECT  0.825 0.525 0.925 0.855 ;
        RECT  0.770 2.540 0.925 3.095 ;
        RECT  0.770 0.525 0.825 1.845 ;
        RECT  0.665 0.525 0.770 3.095 ;
        RECT  0.610 1.685 0.665 2.700 ;
    END
END TLATNCAX4

MACRO TLATNCAX3
    CLASS CORE ;
    FOREIGN TLATNCAX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.345 0.695 5.395 0.945 ;
        RECT  5.245 0.495 5.345 1.125 ;
        RECT  5.085 0.495 5.245 1.860 ;
        RECT  5.035 1.700 5.085 1.860 ;
        RECT  4.875 1.700 5.035 2.710 ;
        RECT  4.775 1.925 4.875 2.710 ;
        RECT  4.725 1.925 4.775 2.400 ;
        END
        ANTENNADIFFAREA     0.6194 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.355 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.2574 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.575 0.395 2.070 ;
        END
        ANTENNAGATEAREA     0.2158 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 -0.250 5.980 0.250 ;
        RECT  5.595 -0.250 5.855 1.125 ;
        RECT  4.785 -0.250 5.595 0.250 ;
        RECT  4.625 -0.250 4.785 0.935 ;
        RECT  3.565 -0.250 4.625 0.250 ;
        RECT  3.305 -0.250 3.565 0.405 ;
        RECT  1.865 -0.250 3.305 0.250 ;
        RECT  1.605 -0.250 1.865 0.755 ;
        RECT  0.385 -0.250 1.605 0.250 ;
        RECT  0.125 -0.250 0.385 1.280 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 3.440 5.980 3.940 ;
        RECT  5.595 2.400 5.855 3.940 ;
        RECT  3.830 3.440 5.595 3.940 ;
        RECT  3.230 3.285 3.830 3.940 ;
        RECT  1.515 3.440 3.230 3.940 ;
        RECT  1.255 2.825 1.515 3.940 ;
        RECT  0.385 3.440 1.255 3.940 ;
        RECT  0.125 2.905 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.585 1.710 5.685 1.970 ;
        RECT  5.425 1.710 5.585 2.220 ;
        RECT  5.415 2.060 5.425 2.220 ;
        RECT  5.255 2.060 5.415 3.050 ;
        RECT  4.335 2.890 5.255 3.050 ;
        RECT  4.605 1.260 4.865 1.520 ;
        RECT  4.445 1.260 4.605 1.420 ;
        RECT  4.285 0.615 4.445 1.420 ;
        RECT  4.175 1.655 4.335 3.050 ;
        RECT  3.145 0.615 4.285 0.775 ;
        RECT  2.840 2.890 4.175 3.050 ;
        RECT  3.995 0.955 4.095 1.215 ;
        RECT  3.835 0.955 3.995 2.115 ;
        RECT  3.645 1.955 3.835 2.115 ;
        RECT  3.495 1.345 3.655 1.635 ;
        RECT  3.485 1.955 3.645 2.215 ;
        RECT  3.145 1.475 3.495 1.635 ;
        RECT  3.325 1.955 3.485 2.585 ;
        RECT  2.985 0.615 3.145 2.425 ;
        RECT  2.685 0.615 2.985 0.775 ;
        RECT  2.495 2.265 2.985 2.425 ;
        RECT  2.680 2.890 2.840 3.220 ;
        RECT  2.645 1.005 2.805 2.085 ;
        RECT  2.425 0.495 2.685 0.775 ;
        RECT  2.055 3.060 2.680 3.220 ;
        RECT  1.325 1.005 2.645 1.165 ;
        RECT  2.545 1.825 2.645 2.085 ;
        RECT  2.235 2.265 2.495 2.865 ;
        RECT  2.305 1.345 2.465 1.605 ;
        RECT  2.055 1.445 2.305 1.605 ;
        RECT  1.895 1.445 2.055 3.220 ;
        RECT  0.895 2.485 1.895 2.645 ;
        RECT  1.295 0.565 1.325 2.195 ;
        RECT  1.175 0.515 1.295 2.195 ;
        RECT  1.165 0.515 1.175 2.295 ;
        RECT  1.035 0.515 1.165 0.775 ;
        RECT  0.915 2.035 1.165 2.295 ;
        RECT  0.825 1.030 0.985 1.660 ;
        RECT  0.735 2.485 0.895 3.165 ;
        RECT  0.665 1.030 0.825 1.290 ;
        RECT  0.735 1.500 0.825 1.660 ;
        RECT  0.635 1.500 0.735 3.165 ;
        RECT  0.575 1.500 0.635 2.645 ;
    END
END TLATNCAX3

MACRO TLATNCAX2
    CLASS CORE ;
    FOREIGN TLATNCAX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.675 2.030 4.935 3.120 ;
        RECT  4.560 2.030 4.675 2.190 ;
        RECT  4.400 0.970 4.560 2.190 ;
        RECT  4.195 0.970 4.400 1.230 ;
        END
        ANTENNADIFFAREA     0.6062 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.355 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.2106 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.575 0.345 2.145 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 -0.250 5.060 0.250 ;
        RECT  4.675 -0.250 4.935 0.405 ;
        RECT  3.915 -0.250 4.675 0.250 ;
        RECT  3.195 -0.250 3.915 0.405 ;
        RECT  1.755 -0.250 3.195 0.250 ;
        RECT  1.495 -0.250 1.755 0.755 ;
        RECT  0.385 -0.250 1.495 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 3.440 5.060 3.940 ;
        RECT  3.815 3.285 4.075 3.940 ;
        RECT  3.310 3.440 3.815 3.940 ;
        RECT  3.050 3.285 3.310 3.940 ;
        RECT  1.470 3.440 3.050 3.940 ;
        RECT  1.210 2.825 1.470 3.940 ;
        RECT  0.385 3.440 1.210 3.940 ;
        RECT  0.125 2.905 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.740 0.595 4.900 1.735 ;
        RECT  3.035 0.595 4.740 0.755 ;
        RECT  4.060 1.465 4.220 2.925 ;
        RECT  2.830 2.765 4.060 2.925 ;
        RECT  3.720 1.135 3.880 2.115 ;
        RECT  3.475 1.135 3.720 1.295 ;
        RECT  3.590 1.955 3.720 2.115 ;
        RECT  3.375 1.955 3.590 2.215 ;
        RECT  3.380 1.480 3.540 1.745 ;
        RECT  3.215 1.035 3.475 1.295 ;
        RECT  3.035 1.585 3.380 1.745 ;
        RECT  3.215 1.955 3.375 2.585 ;
        RECT  2.875 0.595 3.035 2.525 ;
        RECT  2.575 0.595 2.875 0.755 ;
        RECT  2.420 2.365 2.875 2.525 ;
        RECT  2.670 2.765 2.830 3.220 ;
        RECT  2.535 0.935 2.695 2.015 ;
        RECT  1.915 3.060 2.670 3.220 ;
        RECT  2.315 0.495 2.575 0.755 ;
        RECT  1.325 0.935 2.535 1.095 ;
        RECT  2.260 2.365 2.420 2.850 ;
        RECT  2.195 1.275 2.355 1.550 ;
        RECT  2.100 2.690 2.260 2.850 ;
        RECT  2.055 1.390 2.195 1.550 ;
        RECT  1.915 1.390 2.055 2.505 ;
        RECT  1.895 1.390 1.915 3.220 ;
        RECT  1.755 2.345 1.895 3.220 ;
        RECT  1.745 2.345 1.755 2.645 ;
        RECT  0.895 2.485 1.745 2.645 ;
        RECT  1.185 0.935 1.325 2.110 ;
        RECT  1.165 0.495 1.185 2.110 ;
        RECT  1.025 0.495 1.165 1.095 ;
        RECT  1.025 1.950 1.165 2.110 ;
        RECT  0.925 0.495 1.025 0.755 ;
        RECT  0.865 1.950 1.025 2.235 ;
        RECT  0.785 1.470 0.985 1.735 ;
        RECT  0.685 2.485 0.895 3.165 ;
        RECT  0.685 1.005 0.785 1.735 ;
        RECT  0.635 1.005 0.685 3.165 ;
        RECT  0.525 1.005 0.635 2.645 ;
    END
END TLATNCAX2

MACRO CLKMX2X12
    CLASS CORE ;
    FOREIGN CLKMX2X12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.685 1.925 7.695 2.585 ;
        RECT  7.425 1.700 7.685 2.915 ;
        RECT  7.345 1.700 7.425 2.400 ;
        RECT  7.085 0.600 7.345 2.400 ;
        RECT  7.025 1.105 7.085 2.400 ;
        RECT  6.665 1.700 7.025 2.400 ;
        RECT  6.405 1.700 6.665 3.055 ;
        RECT  6.315 1.700 6.405 2.715 ;
        RECT  6.235 1.105 6.315 2.715 ;
        RECT  5.985 0.600 6.235 2.715 ;
        RECT  5.975 0.600 5.985 1.510 ;
        RECT  5.830 2.110 5.985 2.715 ;
        RECT  5.645 2.115 5.830 2.715 ;
        RECT  5.385 2.115 5.645 3.055 ;
        END
        ANTENNADIFFAREA     1.9632 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.585 0.375 2.085 ;
        END
        ANTENNAGATEAREA     0.2457 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 2.925 1.420 3.215 ;
        RECT  1.170 2.925 1.255 3.220 ;
        RECT  1.010 2.925 1.170 3.255 ;
        END
        ANTENNAGATEAREA     0.1703 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 1.480 3.095 1.990 ;
        RECT  2.815 1.315 2.975 1.990 ;
        RECT  2.785 1.480 2.815 1.990 ;
        END
        ANTENNAGATEAREA     0.1703 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.885 -0.250 8.280 0.250 ;
        RECT  7.625 -0.250 7.885 1.170 ;
        RECT  6.795 -0.250 7.625 0.250 ;
        RECT  6.535 -0.250 6.795 1.140 ;
        RECT  5.620 -0.250 6.535 0.250 ;
        RECT  5.360 -0.250 5.620 1.170 ;
        RECT  4.620 -0.250 5.360 0.250 ;
        RECT  4.360 -0.250 4.620 0.405 ;
        RECT  3.420 -0.250 4.360 0.250 ;
        RECT  3.160 -0.250 3.420 1.145 ;
        RECT  0.955 -0.250 3.160 0.250 ;
        RECT  0.695 -0.250 0.955 1.065 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.085 3.440 8.280 3.940 ;
        RECT  7.825 3.285 8.085 3.940 ;
        RECT  7.175 3.440 7.825 3.940 ;
        RECT  6.915 2.615 7.175 3.940 ;
        RECT  6.155 3.440 6.915 3.940 ;
        RECT  5.895 2.930 6.155 3.940 ;
        RECT  5.105 3.440 5.895 3.940 ;
        RECT  4.845 3.285 5.105 3.940 ;
        RECT  4.130 3.440 4.845 3.940 ;
        RECT  3.870 3.285 4.130 3.940 ;
        RECT  2.780 3.440 3.870 3.940 ;
        RECT  2.520 3.285 2.780 3.940 ;
        RECT  0.810 3.440 2.520 3.940 ;
        RECT  0.550 2.930 0.810 3.940 ;
        RECT  0.000 3.440 0.550 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.415 1.575 5.675 1.835 ;
        RECT  5.020 1.575 5.415 1.735 ;
        RECT  4.860 0.865 5.020 2.115 ;
        RECT  4.760 0.865 4.860 1.125 ;
        RECT  4.680 1.955 4.860 2.115 ;
        RECT  4.420 1.955 4.680 2.895 ;
        RECT  3.730 2.735 4.420 2.895 ;
        RECT  4.110 1.535 4.240 1.795 ;
        RECT  3.850 1.035 4.110 1.795 ;
        RECT  3.435 1.635 3.850 1.795 ;
        RECT  3.470 2.705 3.730 2.895 ;
        RECT  3.180 3.085 3.590 3.245 ;
        RECT  3.275 1.635 3.435 2.330 ;
        RECT  3.070 2.170 3.275 2.330 ;
        RECT  3.020 2.945 3.180 3.245 ;
        RECT  1.870 2.945 3.020 3.105 ;
        RECT  2.605 0.845 2.855 1.005 ;
        RECT  2.445 0.845 2.605 2.695 ;
        RECT  2.255 0.435 2.515 0.595 ;
        RECT  2.120 2.535 2.445 2.695 ;
        RECT  2.105 0.930 2.265 2.350 ;
        RECT  2.095 0.435 2.255 0.700 ;
        RECT  1.870 2.190 2.105 2.350 ;
        RECT  1.295 0.540 2.095 0.700 ;
        RECT  1.765 1.065 1.925 2.005 ;
        RECT  1.710 2.190 1.870 3.105 ;
        RECT  1.475 1.065 1.765 1.225 ;
        RECT  1.360 1.845 1.765 2.005 ;
        RECT  1.610 2.190 1.710 2.790 ;
        RECT  1.425 1.405 1.585 1.665 ;
        RECT  1.295 1.405 1.425 1.565 ;
        RECT  1.100 1.845 1.360 2.555 ;
        RECT  1.135 0.540 1.295 1.565 ;
        RECT  0.770 1.245 1.135 1.405 ;
        RECT  0.610 1.245 0.770 2.425 ;
        RECT  0.385 1.245 0.610 1.405 ;
        RECT  0.410 2.265 0.610 2.425 ;
        RECT  0.150 2.265 0.410 2.525 ;
        RECT  0.125 1.015 0.385 1.405 ;
    END
END CLKMX2X12

MACRO CLKMX2X8
    CLASS CORE ;
    FOREIGN CLKMX2X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.290 1.290 6.315 1.990 ;
        RECT  6.230 1.290 6.290 2.345 ;
        RECT  5.970 1.290 6.230 3.055 ;
        RECT  5.855 1.290 5.970 2.400 ;
        RECT  5.850 0.695 5.855 2.400 ;
        RECT  5.830 0.670 5.850 2.400 ;
        RECT  5.590 0.670 5.830 2.345 ;
        RECT  5.210 1.940 5.590 2.345 ;
        RECT  4.950 1.940 5.210 3.055 ;
        END
        ANTENNADIFFAREA     1.3211 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.585 0.375 2.085 ;
        END
        ANTENNAGATEAREA     0.1911 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.150 2.820 1.370 3.220 ;
        RECT  1.045 2.770 1.150 3.220 ;
        RECT  0.990 2.770 1.045 3.030 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.945 1.480 3.095 1.990 ;
        RECT  2.785 1.385 2.945 1.990 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 -0.250 6.900 0.250 ;
        RECT  6.230 -0.250 6.490 0.965 ;
        RECT  5.235 -0.250 6.230 0.250 ;
        RECT  4.975 -0.250 5.235 1.170 ;
        RECT  3.530 -0.250 4.975 0.250 ;
        RECT  3.270 -0.250 3.530 1.145 ;
        RECT  0.955 -0.250 3.270 0.250 ;
        RECT  0.695 -0.250 0.955 1.065 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.740 3.440 6.900 3.940 ;
        RECT  6.480 2.255 6.740 3.940 ;
        RECT  5.720 3.440 6.480 3.940 ;
        RECT  5.460 2.595 5.720 3.940 ;
        RECT  4.670 3.440 5.460 3.940 ;
        RECT  4.410 3.285 4.670 3.940 ;
        RECT  3.695 3.440 4.410 3.940 ;
        RECT  3.435 3.285 3.695 3.940 ;
        RECT  2.785 3.440 3.435 3.940 ;
        RECT  2.525 3.285 2.785 3.940 ;
        RECT  0.810 3.440 2.525 3.940 ;
        RECT  0.550 2.930 0.810 3.940 ;
        RECT  0.000 3.440 0.550 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.635 1.600 5.295 1.760 ;
        RECT  4.630 1.600 4.635 2.140 ;
        RECT  4.470 0.650 4.630 2.140 ;
        RECT  4.370 0.650 4.470 1.250 ;
        RECT  4.245 1.975 4.470 2.140 ;
        RECT  3.985 1.975 4.245 2.915 ;
        RECT  4.110 1.535 4.215 1.795 ;
        RECT  3.860 1.035 4.110 1.795 ;
        RECT  3.850 1.035 3.860 1.295 ;
        RECT  3.445 1.635 3.860 1.795 ;
        RECT  3.335 1.635 3.445 2.520 ;
        RECT  3.285 1.635 3.335 2.600 ;
        RECT  3.075 2.340 3.285 2.600 ;
        RECT  3.010 2.945 3.170 3.240 ;
        RECT  1.920 2.945 3.010 3.105 ;
        RECT  2.695 0.745 2.955 1.075 ;
        RECT  2.605 0.915 2.695 1.075 ;
        RECT  2.445 0.915 2.605 2.695 ;
        RECT  1.295 0.495 2.515 0.655 ;
        RECT  2.120 2.535 2.445 2.695 ;
        RECT  2.105 0.930 2.265 2.350 ;
        RECT  1.920 2.190 2.105 2.350 ;
        RECT  1.765 1.065 1.925 2.005 ;
        RECT  1.760 2.190 1.920 3.105 ;
        RECT  1.735 1.065 1.765 1.225 ;
        RECT  1.360 1.845 1.765 2.005 ;
        RECT  1.610 2.190 1.760 2.450 ;
        RECT  1.475 0.965 1.735 1.225 ;
        RECT  1.425 1.405 1.585 1.665 ;
        RECT  1.295 1.405 1.425 1.565 ;
        RECT  1.100 1.845 1.360 2.555 ;
        RECT  1.135 0.495 1.295 1.565 ;
        RECT  0.770 1.245 1.135 1.405 ;
        RECT  0.610 1.245 0.770 2.425 ;
        RECT  0.385 1.245 0.610 1.405 ;
        RECT  0.410 2.265 0.610 2.425 ;
        RECT  0.150 2.265 0.410 2.525 ;
        RECT  0.125 1.015 0.385 1.405 ;
    END
END CLKMX2X8

MACRO CLKMX2X6
    CLASS CORE ;
    FOREIGN CLKMX2X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.895 1.325 8.155 2.895 ;
        RECT  7.485 1.325 7.895 2.635 ;
        RECT  7.415 1.325 7.485 1.700 ;
        RECT  7.065 2.205 7.485 2.635 ;
        RECT  7.095 0.590 7.415 1.700 ;
        RECT  6.805 2.205 7.065 3.145 ;
        END
        ANTENNADIFFAREA     1.1762 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.590 0.525 1.750 ;
        RECT  0.265 1.590 0.475 1.990 ;
        RECT  0.125 1.700 0.265 1.990 ;
        END
        ANTENNAGATEAREA     0.7124 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.065 1.625 1.485 1.990 ;
        RECT  1.045 1.700 1.065 1.990 ;
        END
        ANTENNAGATEAREA     0.5291 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.085 1.145 6.355 1.660 ;
        END
        ANTENNAGATEAREA     0.5044 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.895 -0.250 8.280 0.250 ;
        RECT  7.635 -0.250 7.895 1.140 ;
        RECT  6.815 -0.250 7.635 0.250 ;
        RECT  6.555 -0.250 6.815 1.140 ;
        RECT  5.725 -0.250 6.555 0.250 ;
        RECT  5.465 -0.250 5.725 0.405 ;
        RECT  1.460 -0.250 5.465 0.250 ;
        RECT  0.860 -0.250 1.460 0.745 ;
        RECT  0.000 -0.250 0.860 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.615 3.440 8.280 3.940 ;
        RECT  7.355 2.865 7.615 3.940 ;
        RECT  6.525 3.440 7.355 3.940 ;
        RECT  6.265 2.935 6.525 3.940 ;
        RECT  5.445 3.440 6.265 3.940 ;
        RECT  5.185 2.955 5.445 3.940 ;
        RECT  1.955 3.440 5.185 3.940 ;
        RECT  1.695 2.555 1.955 3.940 ;
        RECT  0.925 3.440 1.695 3.940 ;
        RECT  0.905 3.285 0.925 3.940 ;
        RECT  0.665 2.640 0.905 3.940 ;
        RECT  0.645 2.640 0.665 2.900 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.815 1.520 6.915 1.780 ;
        RECT  6.655 1.520 6.815 2.025 ;
        RECT  6.505 1.865 6.655 2.025 ;
        RECT  6.345 1.865 6.505 2.670 ;
        RECT  5.045 2.510 6.345 2.670 ;
        RECT  5.885 0.705 6.265 0.965 ;
        RECT  5.885 2.045 5.985 2.305 ;
        RECT  5.725 0.625 5.885 2.305 ;
        RECT  4.795 0.625 5.725 0.785 ;
        RECT  4.535 2.045 5.725 2.205 ;
        RECT  5.370 0.965 5.530 1.865 ;
        RECT  5.095 0.965 5.370 1.125 ;
        RECT  4.115 1.705 5.370 1.865 ;
        RECT  4.455 1.345 5.185 1.505 ;
        RECT  4.945 2.405 5.045 2.670 ;
        RECT  4.785 2.405 4.945 2.985 ;
        RECT  4.635 0.625 4.795 0.965 ;
        RECT  4.025 2.825 4.785 2.985 ;
        RECT  4.275 2.045 4.535 2.645 ;
        RECT  4.295 0.470 4.455 1.505 ;
        RECT  1.925 0.470 4.295 0.630 ;
        RECT  4.025 0.895 4.115 1.865 ;
        RECT  3.955 0.895 4.025 2.985 ;
        RECT  3.865 1.705 3.955 2.985 ;
        RECT  3.765 2.020 3.865 2.985 ;
        RECT  3.005 2.825 3.765 2.985 ;
        RECT  3.515 0.915 3.655 1.175 ;
        RECT  3.355 0.810 3.515 2.620 ;
        RECT  2.565 0.810 3.355 0.970 ;
        RECT  3.255 2.020 3.355 2.620 ;
        RECT  3.005 1.150 3.115 1.310 ;
        RECT  2.845 1.150 3.005 2.985 ;
        RECT  2.745 2.030 2.845 2.985 ;
        RECT  2.495 0.810 2.565 2.375 ;
        RECT  2.405 0.810 2.495 2.905 ;
        RECT  2.155 1.025 2.405 1.285 ;
        RECT  2.235 2.215 2.405 2.905 ;
        RECT  1.415 2.215 2.235 2.375 ;
        RECT  1.925 1.490 2.225 1.650 ;
        RECT  1.765 0.470 1.925 1.650 ;
        RECT  0.865 1.195 1.765 1.355 ;
        RECT  1.155 2.215 1.415 2.905 ;
        RECT  0.705 1.195 0.865 2.355 ;
        RECT  0.390 1.195 0.705 1.355 ;
        RECT  0.385 2.195 0.705 2.355 ;
        RECT  0.385 1.085 0.390 1.355 ;
        RECT  0.125 1.035 0.385 1.355 ;
        RECT  0.125 2.195 0.385 3.145 ;
    END
END CLKMX2X6

MACRO CLKMX2X4
    CLASS CORE ;
    FOREIGN CLKMX2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.105 4.025 2.820 ;
        RECT  3.865 0.470 4.015 2.820 ;
        RECT  3.805 0.470 3.865 1.295 ;
        RECT  3.450 2.660 3.865 2.820 ;
        RECT  3.800 0.695 3.805 1.295 ;
        RECT  3.290 2.660 3.450 2.920 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 0.500 0.610 0.760 ;
        RECT  0.125 0.470 0.335 0.760 ;
        END
        ANTENNAGATEAREA     0.3601 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.495 0.990 2.070 ;
        END
        ANTENNAGATEAREA     0.2496 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 0.880 3.555 1.170 ;
        RECT  3.330 1.010 3.345 1.170 ;
        RECT  3.170 1.010 3.330 1.545 ;
        RECT  3.030 1.285 3.170 1.545 ;
        END
        ANTENNAGATEAREA     0.2613 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 -0.250 4.140 0.250 ;
        RECT  3.240 -0.250 3.500 0.685 ;
        RECT  0.950 -0.250 3.240 0.250 ;
        RECT  0.790 -0.250 0.950 0.715 ;
        RECT  0.000 -0.250 0.790 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 3.440 4.140 3.940 ;
        RECT  3.750 3.005 4.010 3.940 ;
        RECT  2.990 3.440 3.750 3.940 ;
        RECT  2.730 2.985 2.990 3.940 ;
        RECT  0.840 3.440 2.730 3.940 ;
        RECT  0.580 2.895 0.840 3.940 ;
        RECT  0.000 3.440 0.580 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.510 1.575 3.670 2.430 ;
        RECT  3.030 2.270 3.510 2.430 ;
        RECT  2.870 2.270 3.030 2.805 ;
        RECT  2.665 0.880 2.980 1.040 ;
        RECT  2.025 2.645 2.870 2.805 ;
        RECT  2.450 0.435 2.715 0.675 ;
        RECT  2.505 0.880 2.665 2.465 ;
        RECT  2.205 2.305 2.505 2.465 ;
        RECT  1.980 0.515 2.450 0.675 ;
        RECT  2.160 0.895 2.320 2.125 ;
        RECT  2.025 1.965 2.160 2.125 ;
        RECT  1.925 1.965 2.025 2.805 ;
        RECT  1.820 0.515 1.980 1.785 ;
        RECT  1.865 1.965 1.925 3.215 ;
        RECT  1.665 2.275 1.865 3.215 ;
        RECT  1.290 0.515 1.820 0.675 ;
        RECT  1.670 1.575 1.820 1.785 ;
        RECT  1.510 1.575 1.670 1.835 ;
        RECT  1.480 0.860 1.640 1.395 ;
        RECT  1.330 1.235 1.480 1.395 ;
        RECT  1.330 2.255 1.410 3.195 ;
        RECT  1.170 1.235 1.330 3.195 ;
        RECT  1.130 0.515 1.290 1.055 ;
        RECT  1.150 2.255 1.170 3.195 ;
        RECT  0.980 0.895 1.130 1.055 ;
        RECT  0.820 0.895 0.980 1.100 ;
        RECT  0.285 0.940 0.820 1.100 ;
        RECT  0.285 2.170 0.385 2.430 ;
        RECT  0.125 0.940 0.285 2.430 ;
    END
END CLKMX2X4

MACRO CLKMX2X3
    CLASS CORE ;
    FOREIGN CLKMX2X3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 0.880 4.015 1.170 ;
        RECT  3.805 0.880 3.990 1.295 ;
        RECT  3.630 1.035 3.805 1.295 ;
        RECT  3.565 1.135 3.630 1.295 ;
        RECT  3.405 1.135 3.565 2.555 ;
        END
        ANTENNADIFFAREA     0.5960 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 0.520 0.510 0.835 ;
        RECT  0.125 0.470 0.335 0.835 ;
        END
        ANTENNAGATEAREA     0.3328 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.915 1.585 1.075 1.860 ;
        RECT  0.795 1.700 0.915 1.860 ;
        RECT  0.585 1.700 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.2379 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.585 2.885 1.925 ;
        RECT  2.425 1.585 2.635 1.990 ;
        END
        ANTENNAGATEAREA     0.2379 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.350 -0.250 4.140 0.250 ;
        RECT  3.090 -0.250 3.350 0.795 ;
        RECT  0.955 -0.250 3.090 0.250 ;
        RECT  0.695 -0.250 0.955 1.065 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  2.955 3.285 4.015 3.940 ;
        RECT  0.850 3.440 2.955 3.940 ;
        RECT  0.590 2.895 0.850 3.940 ;
        RECT  0.000 3.440 0.590 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.860 1.570 4.020 2.990 ;
        RECT  3.760 1.570 3.860 1.830 ;
        RECT  2.235 2.830 3.860 2.990 ;
        RECT  3.065 1.130 3.225 2.330 ;
        RECT  2.795 1.130 3.065 1.290 ;
        RECT  2.575 2.170 3.065 2.330 ;
        RECT  2.535 1.030 2.795 1.290 ;
        RECT  2.415 2.170 2.575 2.430 ;
        RECT  1.330 0.470 2.455 0.630 ;
        RECT  2.075 0.810 2.235 2.990 ;
        RECT  1.895 2.385 2.075 2.990 ;
        RECT  1.735 0.900 1.895 2.190 ;
        RECT  1.845 2.385 1.895 2.985 ;
        RECT  1.510 0.900 1.735 1.060 ;
        RECT  1.520 2.030 1.735 2.190 ;
        RECT  1.395 1.245 1.555 1.845 ;
        RECT  1.260 2.030 1.520 2.990 ;
        RECT  1.330 1.245 1.395 1.405 ;
        RECT  1.170 0.470 1.330 1.405 ;
        RECT  0.385 1.245 1.170 1.405 ;
        RECT  0.320 2.170 0.420 2.430 ;
        RECT  0.320 1.035 0.385 1.405 ;
        RECT  0.160 1.035 0.320 2.430 ;
        RECT  0.125 1.035 0.160 1.295 ;
    END
END CLKMX2X3

MACRO CLKMX2X2
    CLASS CORE ;
    FOREIGN CLKMX2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.505 1.105 3.555 2.585 ;
        RECT  3.450 0.960 3.505 2.585 ;
        RECT  3.345 0.960 3.450 2.895 ;
        RECT  3.245 0.960 3.345 1.220 ;
        RECT  3.190 1.955 3.345 2.895 ;
        END
        ANTENNADIFFAREA     0.5916 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 2.520 0.455 2.925 ;
        END
        ANTENNAGATEAREA     0.2561 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.700 1.155 1.925 ;
        RECT  0.585 1.700 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.290 2.670 1.820 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 -0.250 3.680 0.250 ;
        RECT  3.180 -0.250 3.440 0.405 ;
        RECT  0.955 -0.250 3.180 0.250 ;
        RECT  0.695 -0.250 0.955 1.180 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 3.440 3.680 3.940 ;
        RECT  2.680 2.725 2.940 3.940 ;
        RECT  0.895 3.440 2.680 3.940 ;
        RECT  0.635 2.200 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.010 1.510 3.150 1.770 ;
        RECT  2.850 0.585 3.010 2.505 ;
        RECT  2.005 0.585 2.850 0.745 ;
        RECT  2.300 2.345 2.850 2.505 ;
        RECT  2.240 0.950 2.550 1.110 ;
        RECT  2.240 2.005 2.430 2.165 ;
        RECT  2.140 2.345 2.300 2.615 ;
        RECT  2.080 0.950 2.240 2.165 ;
        RECT  1.915 2.455 2.140 2.615 ;
        RECT  1.745 0.585 2.005 0.765 ;
        RECT  1.655 2.455 1.915 2.715 ;
        RECT  1.740 1.020 1.900 2.275 ;
        RECT  1.465 1.020 1.740 1.180 ;
        RECT  1.405 2.115 1.740 2.275 ;
        RECT  1.400 1.360 1.560 1.905 ;
        RECT  1.205 0.920 1.465 1.180 ;
        RECT  1.145 2.115 1.405 2.715 ;
        RECT  0.385 1.360 1.400 1.520 ;
        RECT  0.225 0.985 0.385 2.280 ;
        RECT  0.125 0.985 0.225 1.245 ;
        RECT  0.125 2.020 0.225 2.280 ;
    END
END CLKMX2X2

MACRO CLKAND2X12
    CLASS CORE ;
    FOREIGN CLKAND2X12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.315 0.585 5.395 2.585 ;
        RECT  5.055 0.585 5.315 2.735 ;
        RECT  4.755 0.585 5.055 2.055 ;
        RECT  4.495 0.535 4.755 2.055 ;
        RECT  4.295 0.585 4.495 2.055 ;
        RECT  4.265 0.585 4.295 2.735 ;
        RECT  3.675 0.585 4.265 1.145 ;
        RECT  4.035 1.455 4.265 2.735 ;
        RECT  3.415 0.535 3.675 1.145 ;
        RECT  2.315 0.585 3.415 1.145 ;
        END
        ANTENNADIFFAREA     1.8810 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.490 1.605 0.525 1.865 ;
        RECT  0.125 1.605 0.490 2.080 ;
        END
        ANTENNAGATEAREA     0.5642 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 1.705 2.695 1.865 ;
        RECT  1.010 1.290 1.270 1.865 ;
        END
        ANTENNAGATEAREA     0.5642 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.295 -0.250 5.980 0.250 ;
        RECT  5.035 -0.250 5.295 0.405 ;
        RECT  4.215 -0.250 5.035 0.250 ;
        RECT  3.955 -0.250 4.215 0.405 ;
        RECT  3.115 -0.250 3.955 0.250 ;
        RECT  2.855 -0.250 3.115 0.405 ;
        RECT  2.065 -0.250 2.855 0.250 ;
        RECT  1.805 -0.250 2.065 1.085 ;
        RECT  0.385 -0.250 1.805 0.250 ;
        RECT  0.125 -0.250 0.385 1.285 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 3.440 5.980 3.940 ;
        RECT  5.595 2.275 5.855 3.940 ;
        RECT  4.805 3.440 5.595 3.940 ;
        RECT  4.545 2.275 4.805 3.940 ;
        RECT  3.680 3.440 4.545 3.940 ;
        RECT  3.420 1.935 3.680 3.940 ;
        RECT  2.525 3.440 3.420 3.940 ;
        RECT  2.265 2.405 2.525 3.940 ;
        RECT  1.470 3.440 2.265 3.940 ;
        RECT  1.210 2.405 1.470 3.940 ;
        RECT  0.420 3.440 1.210 3.940 ;
        RECT  0.160 2.320 0.420 3.940 ;
        RECT  0.000 3.440 0.160 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.085 1.365 3.525 1.625 ;
        RECT  3.035 1.365 3.085 2.205 ;
        RECT  2.925 1.365 3.035 2.985 ;
        RECT  1.620 1.365 2.925 1.525 ;
        RECT  2.775 2.045 2.925 2.985 ;
        RECT  2.010 2.045 2.775 2.205 ;
        RECT  1.750 2.045 2.010 2.985 ;
        RECT  0.930 2.045 1.750 2.205 ;
        RECT  1.460 0.940 1.620 1.525 ;
        RECT  1.205 0.940 1.460 1.100 ;
        RECT  0.945 0.840 1.205 1.100 ;
        RECT  0.670 2.045 0.930 2.985 ;
    END
END CLKAND2X12

MACRO CLKAND2X8
    CLASS CORE ;
    FOREIGN CLKAND2X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.755 0.585 4.015 2.920 ;
        RECT  3.475 0.585 3.755 2.075 ;
        RECT  3.345 0.535 3.475 2.075 ;
        RECT  3.215 0.535 3.345 0.985 ;
        RECT  2.995 1.675 3.345 2.075 ;
        RECT  2.395 0.585 3.215 0.985 ;
        RECT  2.735 1.675 2.995 3.005 ;
        RECT  2.135 0.535 2.395 0.985 ;
        END
        ANTENNADIFFAREA     1.4004 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.455 1.370 1.615 2.010 ;
        RECT  0.555 1.850 1.455 2.010 ;
        RECT  0.295 1.585 0.555 2.010 ;
        RECT  0.125 1.700 0.295 2.010 ;
        END
        ANTENNAGATEAREA     0.3614 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.290 1.255 1.670 ;
        RECT  0.805 1.410 1.045 1.670 ;
        END
        ANTENNAGATEAREA     0.3614 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 -0.250 4.140 0.250 ;
        RECT  3.755 -0.250 4.015 0.405 ;
        RECT  2.935 -0.250 3.755 0.250 ;
        RECT  2.675 -0.250 2.935 0.405 ;
        RECT  1.885 -0.250 2.675 0.250 ;
        RECT  1.625 -0.250 1.885 0.760 ;
        RECT  0.385 -0.250 1.625 0.250 ;
        RECT  0.125 -0.250 0.385 1.150 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.505 3.440 4.140 3.940 ;
        RECT  3.245 2.255 3.505 3.940 ;
        RECT  2.455 3.440 3.245 3.940 ;
        RECT  2.195 1.725 2.455 3.940 ;
        RECT  1.405 3.440 2.195 3.940 ;
        RECT  1.145 2.635 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.355 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.955 1.165 3.115 1.425 ;
        RECT  1.915 0.950 1.955 2.405 ;
        RECT  1.795 0.950 1.915 2.845 ;
        RECT  1.205 0.950 1.795 1.110 ;
        RECT  1.655 2.245 1.795 2.845 ;
        RECT  0.895 2.245 1.655 2.405 ;
        RECT  0.945 0.850 1.205 1.110 ;
        RECT  0.635 2.245 0.895 2.845 ;
    END
END CLKAND2X8

MACRO CLKAND2X6
    CLASS CORE ;
    FOREIGN CLKAND2X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.055 2.335 3.095 2.995 ;
        RECT  2.795 1.980 3.055 3.085 ;
        RECT  2.635 1.980 2.795 2.330 ;
        RECT  1.975 0.995 2.635 2.330 ;
        RECT  1.845 0.995 1.975 2.920 ;
        RECT  1.755 0.690 1.845 2.920 ;
        RECT  1.585 0.690 1.755 1.290 ;
        RECT  1.715 1.980 1.755 2.920 ;
        END
        ANTENNADIFFAREA     1.1762 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 1.035 1.725 ;
        END
        ANTENNAGATEAREA     0.2522 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.405 1.910 ;
        END
        ANTENNAGATEAREA     0.2522 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.385 -0.250 3.220 0.250 ;
        RECT  2.125 -0.250 2.385 0.795 ;
        RECT  1.305 -0.250 2.125 0.250 ;
        RECT  1.045 -0.250 1.305 0.745 ;
        RECT  0.000 -0.250 1.045 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.515 3.440 3.220 3.940 ;
        RECT  2.255 2.540 2.515 3.940 ;
        RECT  1.455 3.440 2.255 3.940 ;
        RECT  1.155 2.540 1.455 3.940 ;
        RECT  0.385 3.440 1.155 3.940 ;
        RECT  0.125 2.240 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.375 1.510 1.545 1.770 ;
        RECT  1.215 0.950 1.375 2.250 ;
        RECT  0.385 0.950 1.215 1.110 ;
        RECT  0.895 2.090 1.215 2.250 ;
        RECT  0.635 2.090 0.895 3.030 ;
        RECT  0.125 0.850 0.385 1.110 ;
    END
END CLKAND2X6

MACRO CLKAND2X4
    CLASS CORE ;
    FOREIGN CLKAND2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.005 0.880 2.175 1.770 ;
        RECT  1.845 0.880 2.005 3.210 ;
        RECT  1.745 0.495 1.845 3.210 ;
        RECT  1.585 0.495 1.745 1.120 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.650 1.095 1.935 ;
        RECT  0.610 1.650 0.795 1.990 ;
        RECT  0.585 1.700 0.610 1.990 ;
        END
        ANTENNAGATEAREA     0.1833 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.545 0.385 2.105 ;
        END
        ANTENNAGATEAREA     0.1833 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.335 -0.250 2.760 0.250 ;
        RECT  1.075 -0.250 1.335 1.115 ;
        RECT  0.000 -0.250 1.075 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 3.440 2.760 3.940 ;
        RECT  2.285 2.215 2.545 3.940 ;
        RECT  1.465 3.440 2.285 3.940 ;
        RECT  1.205 2.610 1.465 3.940 ;
        RECT  0.385 3.440 1.205 3.940 ;
        RECT  0.125 2.445 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.450 1.565 1.530 1.825 ;
        RECT  1.290 1.310 1.450 2.370 ;
        RECT  0.725 1.310 1.290 1.470 ;
        RECT  0.925 2.210 1.290 2.370 ;
        RECT  0.665 2.210 0.925 2.810 ;
        RECT  0.565 1.075 0.725 1.470 ;
        RECT  0.415 1.075 0.565 1.235 ;
        RECT  0.155 0.975 0.415 1.235 ;
    END
END CLKAND2X4

MACRO CLKAND2X3
    CLASS CORE ;
    FOREIGN CLKAND2X3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 0.680 1.865 1.280 ;
        RECT  1.725 0.680 1.765 2.310 ;
        RECT  1.605 0.680 1.725 2.725 ;
        RECT  1.505 2.110 1.605 2.725 ;
        RECT  1.465 2.125 1.505 2.725 ;
        END
        ANTENNADIFFAREA     0.5926 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.825 2.800 0.925 3.060 ;
        RECT  0.795 2.585 0.825 3.060 ;
        RECT  0.665 2.520 0.795 3.060 ;
        RECT  0.585 2.520 0.665 2.810 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.600 0.445 1.860 ;
        RECT  0.125 1.600 0.335 2.265 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.325 -0.250 2.300 0.250 ;
        RECT  1.065 -0.250 1.325 0.885 ;
        RECT  0.000 -0.250 1.065 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 3.440 2.300 3.940 ;
        RECT  1.865 3.285 2.125 3.940 ;
        RECT  1.325 3.440 1.865 3.940 ;
        RECT  1.065 3.285 1.325 3.940 ;
        RECT  0.385 3.440 1.065 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.055 1.590 1.385 1.860 ;
        RECT  0.895 1.130 1.055 2.220 ;
        RECT  0.475 1.130 0.895 1.290 ;
        RECT  0.785 2.060 0.895 2.220 ;
        RECT  0.525 2.060 0.785 2.320 ;
        RECT  0.215 1.030 0.475 1.290 ;
    END
END CLKAND2X3

MACRO CLKAND2X2
    CLASS CORE ;
    FOREIGN CLKAND2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.515 2.175 2.585 ;
        RECT  2.010 1.115 2.100 2.585 ;
        RECT  1.940 1.115 2.010 2.970 ;
        RECT  1.835 1.115 1.940 1.275 ;
        RECT  1.750 2.030 1.940 2.970 ;
        RECT  1.575 1.015 1.835 1.275 ;
        END
        ANTENNADIFFAREA     0.5882 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.735 2.520 1.015 3.035 ;
        RECT  0.585 2.520 0.735 2.810 ;
        END
        ANTENNAGATEAREA     0.0923 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.465 0.430 1.835 ;
        RECT  0.135 1.465 0.335 1.990 ;
        RECT  0.125 1.700 0.135 1.990 ;
        END
        ANTENNAGATEAREA     0.0923 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 -0.250 2.300 0.250 ;
        RECT  1.030 -0.250 1.290 1.135 ;
        RECT  0.000 -0.250 1.030 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 3.440 2.300 3.940 ;
        RECT  1.205 2.030 1.465 3.940 ;
        RECT  0.385 3.440 1.205 3.940 ;
        RECT  0.125 2.170 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.410 1.590 1.670 1.850 ;
        RECT  0.925 1.690 1.410 1.850 ;
        RECT  0.825 1.690 0.925 2.275 ;
        RECT  0.665 1.115 0.825 2.275 ;
        RECT  0.410 1.115 0.665 1.275 ;
        RECT  0.150 1.015 0.410 1.275 ;
    END
END CLKAND2X2

MACRO CLKINVX20
    CLASS CORE ;
    FOREIGN CLKINVX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.090 1.105 8.155 2.995 ;
        RECT  7.830 0.865 8.090 3.215 ;
        RECT  7.035 0.865 7.830 1.990 ;
        RECT  6.775 0.865 7.035 3.215 ;
        RECT  6.015 0.865 6.775 1.990 ;
        RECT  5.755 0.865 6.015 2.935 ;
        RECT  5.200 0.865 5.755 2.770 ;
        RECT  5.185 0.645 5.200 2.770 ;
        RECT  4.940 0.645 5.185 1.405 ;
        RECT  4.995 2.170 5.185 2.770 ;
        RECT  4.735 2.170 4.995 3.215 ;
        RECT  4.180 0.865 4.940 1.405 ;
        RECT  4.725 2.170 4.735 2.995 ;
        RECT  4.015 2.170 4.725 2.770 ;
        RECT  3.920 0.645 4.180 1.405 ;
        RECT  3.975 2.170 4.015 2.995 ;
        RECT  3.715 2.170 3.975 3.215 ;
        RECT  3.160 0.865 3.920 1.405 ;
        RECT  2.950 2.170 3.715 2.770 ;
        RECT  2.900 0.645 3.160 1.405 ;
        RECT  2.690 2.170 2.950 3.195 ;
        RECT  2.885 0.695 2.900 1.405 ;
        RECT  2.110 0.865 2.885 1.405 ;
        RECT  1.920 2.170 2.690 2.770 ;
        RECT  1.850 0.645 2.110 1.405 ;
        RECT  1.660 2.170 1.920 3.195 ;
        RECT  1.090 0.865 1.850 1.405 ;
        RECT  0.640 2.170 1.660 2.770 ;
        RECT  0.830 0.685 1.090 1.405 ;
        RECT  0.585 2.335 0.640 2.585 ;
        END
        ANTENNADIFFAREA     6.3195 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.630 4.845 1.790 ;
        RECT  3.345 1.630 3.555 1.990 ;
        RECT  0.845 1.630 3.345 1.790 ;
        END
        ANTENNAGATEAREA     4.2042 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.710 -0.250 8.740 0.250 ;
        RECT  5.450 -0.250 5.710 0.685 ;
        RECT  4.690 -0.250 5.450 0.250 ;
        RECT  4.430 -0.250 4.690 0.685 ;
        RECT  3.670 -0.250 4.430 0.250 ;
        RECT  3.410 -0.250 3.670 0.685 ;
        RECT  2.620 -0.250 3.410 0.250 ;
        RECT  2.360 -0.250 2.620 0.685 ;
        RECT  1.600 -0.250 2.360 0.250 ;
        RECT  1.340 -0.250 1.600 0.685 ;
        RECT  0.580 -0.250 1.340 0.250 ;
        RECT  0.320 -0.250 0.580 1.275 ;
        RECT  0.000 -0.250 0.320 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.600 3.440 8.740 3.940 ;
        RECT  8.340 2.275 8.600 3.940 ;
        RECT  7.575 3.440 8.340 3.940 ;
        RECT  7.315 2.275 7.575 3.940 ;
        RECT  6.525 3.440 7.315 3.940 ;
        RECT  6.265 2.275 6.525 3.940 ;
        RECT  5.505 3.440 6.265 3.940 ;
        RECT  5.245 2.950 5.505 3.940 ;
        RECT  4.485 3.440 5.245 3.940 ;
        RECT  4.225 2.950 4.485 3.940 ;
        RECT  3.460 3.440 4.225 3.940 ;
        RECT  3.200 2.950 3.460 3.940 ;
        RECT  2.440 3.440 3.200 3.940 ;
        RECT  2.180 2.950 2.440 3.940 ;
        RECT  1.410 3.440 2.180 3.940 ;
        RECT  1.150 2.950 1.410 3.940 ;
        RECT  0.390 3.440 1.150 3.940 ;
        RECT  0.130 2.195 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
END CLKINVX20

MACRO CLKINVX16
    CLASS CORE ;
    FOREIGN CLKINVX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.065 1.105 7.235 2.995 ;
        RECT  6.805 0.865 7.065 3.215 ;
        RECT  6.010 0.865 6.805 2.020 ;
        RECT  5.750 0.865 6.010 3.215 ;
        RECT  4.990 0.865 5.750 2.020 ;
        RECT  4.730 0.865 4.990 2.935 ;
        RECT  4.175 0.865 4.730 2.770 ;
        RECT  4.165 0.645 4.175 2.770 ;
        RECT  3.915 0.645 4.165 1.405 ;
        RECT  4.015 2.110 4.165 2.770 ;
        RECT  3.990 2.110 4.015 2.995 ;
        RECT  3.970 2.170 3.990 2.995 ;
        RECT  3.710 2.170 3.970 3.215 ;
        RECT  3.155 0.865 3.915 1.405 ;
        RECT  2.950 2.170 3.710 2.770 ;
        RECT  2.895 0.645 3.155 1.405 ;
        RECT  2.690 2.170 2.950 3.215 ;
        RECT  2.885 0.695 2.895 1.405 ;
        RECT  2.135 0.865 2.885 1.405 ;
        RECT  1.925 2.170 2.690 2.770 ;
        RECT  1.875 0.645 2.135 1.405 ;
        RECT  1.665 2.170 1.925 3.195 ;
        RECT  1.085 0.865 1.875 1.405 ;
        RECT  0.895 2.170 1.665 2.770 ;
        RECT  0.825 0.685 1.085 1.405 ;
        RECT  0.635 2.170 0.895 2.835 ;
        RECT  0.585 2.335 0.635 2.585 ;
        END
        ANTENNADIFFAREA     5.2074 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.630 3.945 1.790 ;
        RECT  2.425 1.630 2.635 1.990 ;
        RECT  0.965 1.630 2.425 1.790 ;
        END
        ANTENNAGATEAREA     3.3579 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.685 -0.250 7.360 0.250 ;
        RECT  4.425 -0.250 4.685 0.685 ;
        RECT  3.665 -0.250 4.425 0.250 ;
        RECT  3.405 -0.250 3.665 0.685 ;
        RECT  2.645 -0.250 3.405 0.250 ;
        RECT  2.385 -0.250 2.645 0.685 ;
        RECT  1.595 -0.250 2.385 0.250 ;
        RECT  1.335 -0.250 1.595 0.685 ;
        RECT  0.575 -0.250 1.335 0.250 ;
        RECT  0.315 -0.250 0.575 1.275 ;
        RECT  0.000 -0.250 0.315 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.550 3.440 7.360 3.940 ;
        RECT  6.290 2.275 6.550 3.940 ;
        RECT  5.500 3.440 6.290 3.940 ;
        RECT  5.240 2.275 5.500 3.940 ;
        RECT  4.480 3.440 5.240 3.940 ;
        RECT  4.220 2.950 4.480 3.940 ;
        RECT  3.460 3.440 4.220 3.940 ;
        RECT  3.200 2.950 3.460 3.940 ;
        RECT  2.435 3.440 3.200 3.940 ;
        RECT  2.175 2.950 2.435 3.940 ;
        RECT  1.415 3.440 2.175 3.940 ;
        RECT  1.155 2.950 1.415 3.940 ;
        RECT  0.385 3.440 1.155 3.940 ;
        RECT  0.125 2.265 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END CLKINVX16

MACRO CLKINVX12
    CLASS CORE ;
    FOREIGN CLKINVX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.315 1.105 5.395 2.995 ;
        RECT  5.055 0.865 5.315 3.215 ;
        RECT  4.910 0.865 5.055 1.990 ;
        RECT  4.295 0.865 4.910 1.815 ;
        RECT  4.035 0.865 4.295 2.915 ;
        RECT  3.480 0.865 4.035 2.645 ;
        RECT  3.345 0.645 3.480 2.645 ;
        RECT  3.220 0.645 3.345 1.405 ;
        RECT  3.275 2.170 3.345 2.645 ;
        RECT  3.015 2.170 3.275 3.215 ;
        RECT  2.460 0.865 3.220 1.405 ;
        RECT  2.255 2.170 3.015 2.645 ;
        RECT  2.200 0.645 2.460 1.405 ;
        RECT  1.995 2.170 2.255 3.215 ;
        RECT  1.440 0.865 2.200 1.405 ;
        RECT  1.965 2.170 1.995 2.995 ;
        RECT  1.230 2.170 1.965 2.645 ;
        RECT  1.180 0.645 1.440 1.405 ;
        RECT  0.970 2.170 1.230 2.835 ;
        END
        ANTENNADIFFAREA     3.7372 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.630 3.100 1.790 ;
        RECT  1.965 1.630 2.175 1.990 ;
        RECT  0.800 1.630 1.965 1.790 ;
        END
        ANTENNAGATEAREA     2.4882 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 -0.250 5.980 0.250 ;
        RECT  3.730 -0.250 3.990 0.685 ;
        RECT  2.970 -0.250 3.730 0.250 ;
        RECT  2.710 -0.250 2.970 0.685 ;
        RECT  1.950 -0.250 2.710 0.250 ;
        RECT  1.690 -0.250 1.950 0.685 ;
        RECT  0.900 -0.250 1.690 0.250 ;
        RECT  0.640 -0.250 0.900 1.135 ;
        RECT  0.000 -0.250 0.640 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 3.440 5.980 3.940 ;
        RECT  5.595 2.275 5.855 3.940 ;
        RECT  4.805 3.440 5.595 3.940 ;
        RECT  4.545 2.275 4.805 3.940 ;
        RECT  3.785 3.440 4.545 3.940 ;
        RECT  3.525 2.950 3.785 3.940 ;
        RECT  2.765 3.440 3.525 3.940 ;
        RECT  2.505 2.950 2.765 3.940 ;
        RECT  1.740 3.440 2.505 3.940 ;
        RECT  1.480 2.950 1.740 3.940 ;
        RECT  0.720 3.440 1.480 3.940 ;
        RECT  0.460 2.075 0.720 3.940 ;
        RECT  0.000 3.440 0.460 3.940 ;
        END
    END VDD
END CLKINVX12

MACRO CLKINVX8
    CLASS CORE ;
    FOREIGN CLKINVX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.290 2.635 1.990 ;
        RECT  2.155 0.695 2.175 2.175 ;
        RECT  1.995 0.685 2.155 2.465 ;
        RECT  1.855 0.685 1.995 3.005 ;
        RECT  1.725 0.965 1.855 3.005 ;
        RECT  1.720 0.965 1.725 1.720 ;
        RECT  1.695 2.065 1.725 3.005 ;
        RECT  1.015 0.965 1.720 1.365 ;
        RECT  0.915 2.065 1.695 2.465 ;
        RECT  0.715 0.685 1.015 1.365 ;
        RECT  0.615 2.065 0.915 3.020 ;
        RECT  0.585 2.335 0.615 2.585 ;
        END
        ANTENNADIFFAREA     1.4828 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 1.585 1.510 1.845 ;
        RECT  0.335 1.585 0.385 1.975 ;
        RECT  0.125 1.585 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.8996 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 -0.250 2.760 0.250 ;
        RECT  1.305 -0.250 1.565 0.745 ;
        RECT  0.425 -0.250 1.305 0.250 ;
        RECT  0.165 -0.250 0.425 1.160 ;
        RECT  0.000 -0.250 0.165 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.515 3.440 2.760 3.940 ;
        RECT  2.255 2.765 2.515 3.940 ;
        RECT  1.435 3.440 2.255 3.940 ;
        RECT  1.175 2.725 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.255 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END CLKINVX8

MACRO CLKINVX6
    CLASS CORE ;
    FOREIGN CLKINVX6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.105 2.175 2.585 ;
        RECT  1.790 0.905 2.150 2.895 ;
        RECT  1.095 1.005 1.790 2.305 ;
        RECT  1.085 0.905 1.095 2.305 ;
        RECT  1.045 0.905 1.085 2.895 ;
        RECT  0.735 0.905 1.045 1.365 ;
        RECT  0.725 1.945 1.045 2.895 ;
        END
        ANTENNADIFFAREA     1.2456 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.575 0.865 1.735 ;
        RECT  0.175 1.290 0.335 1.735 ;
        RECT  0.125 1.290 0.175 1.580 ;
        END
        ANTENNAGATEAREA     0.6747 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 -0.250 2.300 0.250 ;
        RECT  1.315 -0.250 1.575 0.795 ;
        RECT  0.495 -0.250 1.315 0.250 ;
        RECT  0.235 -0.250 0.495 0.815 ;
        RECT  0.000 -0.250 0.235 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 3.440 2.300 3.940 ;
        RECT  1.315 2.525 1.575 3.940 ;
        RECT  0.495 3.440 1.315 3.940 ;
        RECT  0.235 2.200 0.495 3.940 ;
        RECT  0.000 3.440 0.235 3.940 ;
        END
    END VDD
END CLKINVX6

MACRO CLKINVX4
    CLASS CORE ;
    FOREIGN CLKINVX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.115 0.880 1.265 2.035 ;
        RECT  1.025 0.640 1.115 2.035 ;
        RECT  0.855 0.640 1.025 1.240 ;
        RECT  0.965 1.795 1.025 2.035 ;
        RECT  0.705 1.795 0.965 2.910 ;
        END
        ANTENNADIFFAREA     0.7804 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.455 0.845 1.615 ;
        RECT  0.175 1.455 0.335 1.990 ;
        RECT  0.125 1.700 0.175 1.990 ;
        END
        ANTENNAGATEAREA     0.4420 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.570 -0.250 1.840 0.250 ;
        RECT  0.310 -0.250 0.570 1.170 ;
        RECT  0.000 -0.250 0.310 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 3.440 1.840 3.940 ;
        RECT  1.245 2.215 1.505 3.940 ;
        RECT  0.425 3.440 1.245 3.940 ;
        RECT  0.165 2.210 0.425 3.940 ;
        RECT  0.000 3.440 0.165 3.940 ;
        END
    END VDD
END CLKINVX4

MACRO CLKINVX3
    CLASS CORE ;
    FOREIGN CLKINVX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.380 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.700 1.255 1.990 ;
        RECT  0.820 0.695 0.980 2.365 ;
        RECT  0.720 0.695 0.820 1.295 ;
        RECT  0.770 2.110 0.820 2.805 ;
        RECT  0.560 2.205 0.770 2.805 ;
        END
        ANTENNADIFFAREA     0.5892 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.355 1.600 0.615 1.860 ;
        RECT  0.335 1.700 0.355 1.860 ;
        RECT  0.125 1.700 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.3354 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.425 -0.250 1.380 0.250 ;
        RECT  0.165 -0.250 0.425 1.175 ;
        RECT  0.000 -0.250 0.165 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 3.440 1.380 3.940 ;
        RECT  0.995 3.285 1.255 3.940 ;
        RECT  0.385 3.440 0.995 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END CLKINVX3

MACRO CLKINVX2
    CLASS CORE ;
    FOREIGN CLKINVX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.380 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.050 1.700 1.255 1.990 ;
        RECT  0.890 1.035 1.050 2.895 ;
        RECT  0.790 1.035 0.890 1.295 ;
        RECT  0.790 1.955 0.890 2.895 ;
        END
        ANTENNADIFFAREA     0.5882 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.585 0.595 1.845 ;
        RECT  0.125 1.585 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 -0.250 1.380 0.250 ;
        RECT  0.250 -0.250 0.510 1.190 ;
        RECT  0.000 -0.250 0.250 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 3.440 1.380 3.940 ;
        RECT  0.250 2.190 0.510 3.940 ;
        RECT  0.000 3.440 0.250 3.940 ;
        END
    END VDD
END CLKINVX2

MACRO CLKINVX1
    CLASS CORE ;
    FOREIGN CLKINVX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 0.775 0.795 2.680 ;
        RECT  0.535 0.775 0.585 1.035 ;
        RECT  0.535 2.080 0.585 2.680 ;
        END
        ANTENNADIFFAREA     0.4012 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.405 0.405 1.665 ;
        RECT  0.145 1.405 0.335 1.990 ;
        RECT  0.125 1.515 0.145 1.990 ;
        END
        ANTENNAGATEAREA     0.1534 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.250 0.920 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 0.920 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END CLKINVX1

MACRO CLKBUFX20
    CLASS CORE ;
    FOREIGN CLKBUFX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.340 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.005 1.835 12.955 2.435 ;
        RECT  11.745 1.835 12.005 2.980 ;
        RECT  10.985 1.835 11.745 2.435 ;
        RECT  10.725 1.835 10.985 2.980 ;
        RECT  10.705 1.835 10.725 2.585 ;
        RECT  9.995 1.835 10.705 2.435 ;
        RECT  9.965 1.835 9.995 2.585 ;
        RECT  9.705 1.835 9.965 2.980 ;
        RECT  9.075 1.835 9.705 2.435 ;
        RECT  8.945 1.290 9.075 2.435 ;
        RECT  8.685 1.290 8.945 2.980 ;
        RECT  8.195 1.290 8.685 2.435 ;
        RECT  7.925 0.585 8.195 2.435 ;
        RECT  7.665 0.585 7.925 2.980 ;
        RECT  7.295 0.585 7.665 2.435 ;
        RECT  3.585 0.585 7.295 1.185 ;
        RECT  6.905 1.835 7.295 2.435 ;
        RECT  6.645 1.835 6.905 2.980 ;
        RECT  5.885 1.835 6.645 2.435 ;
        RECT  5.625 1.835 5.885 2.980 ;
        RECT  4.935 1.835 5.625 2.435 ;
        RECT  4.865 1.835 4.935 2.585 ;
        RECT  4.605 1.835 4.865 2.980 ;
        RECT  3.845 1.835 4.605 2.435 ;
        RECT  3.585 1.835 3.845 2.980 ;
        END
        ANTENNADIFFAREA     6.2120 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.495 2.995 1.755 ;
        RECT  0.585 1.290 0.795 1.755 ;
        RECT  0.355 1.495 0.585 1.755 ;
        END
        ANTENNAGATEAREA     1.3104 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.675 -0.250 13.340 0.250 ;
        RECT  8.415 -0.250 8.675 1.095 ;
        RECT  7.625 -0.250 8.415 0.250 ;
        RECT  7.365 -0.250 7.625 0.405 ;
        RECT  6.545 -0.250 7.365 0.250 ;
        RECT  6.285 -0.250 6.545 0.405 ;
        RECT  5.465 -0.250 6.285 0.250 ;
        RECT  5.205 -0.250 5.465 0.405 ;
        RECT  4.385 -0.250 5.205 0.250 ;
        RECT  4.125 -0.250 4.385 0.405 ;
        RECT  3.335 -0.250 4.125 0.250 ;
        RECT  3.075 -0.250 3.335 0.755 ;
        RECT  2.315 -0.250 3.075 0.250 ;
        RECT  2.055 -0.250 2.315 0.740 ;
        RECT  0.000 -0.250 2.055 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.570 3.440 13.340 3.940 ;
        RECT  12.310 2.735 12.570 3.940 ;
        RECT  11.495 3.440 12.310 3.940 ;
        RECT  11.235 2.615 11.495 3.940 ;
        RECT  10.475 3.440 11.235 3.940 ;
        RECT  10.215 2.615 10.475 3.940 ;
        RECT  9.455 3.440 10.215 3.940 ;
        RECT  9.195 2.615 9.455 3.940 ;
        RECT  8.435 3.440 9.195 3.940 ;
        RECT  8.175 2.615 8.435 3.940 ;
        RECT  7.415 3.440 8.175 3.940 ;
        RECT  7.155 2.615 7.415 3.940 ;
        RECT  6.395 3.440 7.155 3.940 ;
        RECT  6.135 2.615 6.395 3.940 ;
        RECT  5.375 3.440 6.135 3.940 ;
        RECT  5.115 2.615 5.375 3.940 ;
        RECT  4.355 3.440 5.115 3.940 ;
        RECT  4.095 2.615 4.355 3.940 ;
        RECT  3.335 3.440 4.095 3.940 ;
        RECT  3.075 2.275 3.335 3.940 ;
        RECT  2.315 3.440 3.075 3.940 ;
        RECT  2.055 2.275 2.315 3.940 ;
        RECT  1.295 3.440 2.055 3.940 ;
        RECT  1.035 2.275 1.295 3.940 ;
        RECT  0.385 3.440 1.035 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.335 1.455 7.075 1.615 ;
        RECT  3.175 1.135 3.335 2.095 ;
        RECT  2.825 1.135 3.175 1.295 ;
        RECT  2.825 1.935 3.175 2.095 ;
        RECT  2.565 0.695 2.825 1.295 ;
        RECT  2.565 1.935 2.825 3.025 ;
        RECT  1.805 1.135 2.565 1.295 ;
        RECT  1.805 1.935 2.565 2.095 ;
        RECT  1.545 0.695 1.805 1.295 ;
        RECT  1.545 1.935 1.805 3.025 ;
        RECT  0.785 1.935 1.545 2.095 ;
        RECT  0.625 1.935 0.785 2.535 ;
        RECT  0.525 2.275 0.625 2.535 ;
    END
END CLKBUFX20

MACRO CLKBUFX16
    CLASS CORE ;
    FOREIGN CLKBUFX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 1.835 9.565 2.895 ;
        RECT  8.615 1.835 9.305 2.435 ;
        RECT  8.545 1.835 8.615 2.585 ;
        RECT  8.285 1.835 8.545 2.895 ;
        RECT  7.525 1.835 8.285 2.435 ;
        RECT  7.265 1.835 7.525 2.895 ;
        RECT  7.235 1.835 7.265 2.435 ;
        RECT  6.685 1.290 7.235 2.435 ;
        RECT  6.505 0.585 6.685 2.435 ;
        RECT  6.245 0.585 6.505 2.895 ;
        RECT  6.105 0.585 6.245 2.435 ;
        RECT  3.185 0.585 6.105 1.185 ;
        RECT  5.485 1.835 6.105 2.435 ;
        RECT  5.225 1.835 5.485 2.895 ;
        RECT  5.185 1.835 5.225 2.585 ;
        RECT  4.475 1.835 5.185 2.435 ;
        RECT  4.465 1.835 4.475 2.585 ;
        RECT  4.205 1.835 4.465 2.895 ;
        RECT  3.445 1.835 4.205 2.435 ;
        RECT  3.185 1.835 3.445 2.895 ;
        END
        ANTENNADIFFAREA     4.7348 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.495 2.425 1.755 ;
        RECT  0.585 1.290 0.795 1.755 ;
        RECT  0.465 1.495 0.585 1.755 ;
        END
        ANTENNAGATEAREA     1.0556 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.195 -0.250 10.580 0.250 ;
        RECT  6.935 -0.250 7.195 1.095 ;
        RECT  6.145 -0.250 6.935 0.250 ;
        RECT  5.885 -0.250 6.145 0.405 ;
        RECT  5.065 -0.250 5.885 0.250 ;
        RECT  4.805 -0.250 5.065 0.405 ;
        RECT  3.985 -0.250 4.805 0.250 ;
        RECT  3.725 -0.250 3.985 0.405 ;
        RECT  2.935 -0.250 3.725 0.250 ;
        RECT  2.675 -0.250 2.935 0.775 ;
        RECT  1.915 -0.250 2.675 0.250 ;
        RECT  1.655 -0.250 1.915 0.975 ;
        RECT  0.000 -0.250 1.655 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.075 3.440 10.580 3.940 ;
        RECT  9.815 2.275 10.075 3.940 ;
        RECT  9.055 3.440 9.815 3.940 ;
        RECT  8.795 2.615 9.055 3.940 ;
        RECT  8.035 3.440 8.795 3.940 ;
        RECT  7.775 2.615 8.035 3.940 ;
        RECT  7.015 3.440 7.775 3.940 ;
        RECT  6.755 2.615 7.015 3.940 ;
        RECT  5.995 3.440 6.755 3.940 ;
        RECT  5.735 2.615 5.995 3.940 ;
        RECT  4.975 3.440 5.735 3.940 ;
        RECT  4.715 2.615 4.975 3.940 ;
        RECT  3.955 3.440 4.715 3.940 ;
        RECT  3.695 2.615 3.955 3.940 ;
        RECT  2.935 3.440 3.695 3.940 ;
        RECT  2.675 2.275 2.935 3.940 ;
        RECT  1.915 3.440 2.675 3.940 ;
        RECT  1.655 2.275 1.915 3.940 ;
        RECT  0.895 3.440 1.655 3.940 ;
        RECT  0.635 2.455 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.765 1.455 5.655 1.615 ;
        RECT  2.605 1.155 2.765 2.095 ;
        RECT  2.425 1.155 2.605 1.315 ;
        RECT  2.425 1.935 2.605 2.095 ;
        RECT  2.165 0.695 2.425 1.315 ;
        RECT  2.165 1.935 2.425 2.980 ;
        RECT  1.405 1.155 2.165 1.315 ;
        RECT  1.405 1.935 2.165 2.095 ;
        RECT  1.245 0.815 1.405 1.315 ;
        RECT  1.145 1.935 1.405 3.130 ;
        RECT  1.145 0.815 1.245 1.075 ;
        RECT  0.385 1.935 1.145 2.095 ;
        RECT  0.125 1.935 0.385 2.555 ;
    END
END CLKBUFX16

MACRO CLKBUFX12
    CLASS CORE ;
    FOREIGN CLKBUFX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.570 1.290 6.775 2.085 ;
        RECT  6.315 0.585 6.570 2.085 ;
        RECT  6.235 0.585 6.315 2.585 ;
        RECT  6.105 0.585 6.235 3.025 ;
        RECT  3.075 0.585 6.105 1.035 ;
        RECT  5.975 1.635 6.105 3.025 ;
        RECT  5.155 1.635 5.975 2.085 ;
        RECT  4.895 1.635 5.155 3.025 ;
        RECT  4.135 1.635 4.895 2.085 ;
        RECT  3.875 1.635 4.135 3.025 ;
        RECT  3.805 1.635 3.875 2.585 ;
        RECT  3.655 1.635 3.805 2.435 ;
        RECT  3.115 1.985 3.655 2.435 ;
        RECT  2.855 1.985 3.115 3.145 ;
        RECT  2.625 0.585 3.075 1.385 ;
        RECT  1.915 0.935 2.625 1.385 ;
        RECT  1.655 0.675 1.915 1.385 ;
        END
        ANTENNADIFFAREA     3.4747 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.520 1.135 1.780 ;
        RECT  0.125 1.290 0.335 1.780 ;
        END
        ANTENNAGATEAREA     0.7800 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 -0.250 6.900 0.250 ;
        RECT  6.515 -0.250 6.775 0.405 ;
        RECT  5.665 -0.250 6.515 0.250 ;
        RECT  5.405 -0.250 5.665 0.405 ;
        RECT  4.555 -0.250 5.405 0.250 ;
        RECT  4.295 -0.250 4.555 0.405 ;
        RECT  3.475 -0.250 4.295 0.250 ;
        RECT  3.215 -0.250 3.475 0.405 ;
        RECT  2.425 -0.250 3.215 0.250 ;
        RECT  2.165 -0.250 2.425 0.755 ;
        RECT  1.405 -0.250 2.165 0.250 ;
        RECT  1.145 -0.250 1.405 0.935 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.110 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.275 6.775 3.940 ;
        RECT  5.695 3.440 6.515 3.940 ;
        RECT  5.435 2.275 5.695 3.940 ;
        RECT  4.645 3.440 5.435 3.940 ;
        RECT  4.385 2.275 4.645 3.940 ;
        RECT  3.625 3.440 4.385 3.940 ;
        RECT  3.365 2.615 3.625 3.940 ;
        RECT  2.515 3.440 3.365 3.940 ;
        RECT  2.255 2.070 2.515 3.940 ;
        RECT  1.405 3.440 2.255 3.940 ;
        RECT  1.145 2.420 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.160 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.435 1.255 5.915 1.415 ;
        RECT  3.275 1.255 3.435 1.765 ;
        RECT  1.475 1.605 3.275 1.765 ;
        RECT  1.655 1.995 1.915 3.020 ;
        RECT  1.475 1.995 1.655 2.155 ;
        RECT  1.315 1.135 1.475 2.155 ;
        RECT  0.895 1.135 1.315 1.295 ;
        RECT  0.895 1.995 1.315 2.155 ;
        RECT  0.635 0.675 0.895 1.295 ;
        RECT  0.635 1.995 0.895 2.935 ;
    END
END CLKBUFX12

MACRO CLKBUFX8
    CLASS CORE ;
    FOREIGN CLKBUFX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.035 1.105 3.095 1.990 ;
        RECT  2.825 0.635 3.035 1.990 ;
        RECT  2.775 0.635 2.825 2.375 ;
        RECT  2.690 0.880 2.775 2.375 ;
        RECT  2.610 0.880 2.690 2.915 ;
        RECT  2.430 0.940 2.610 2.915 ;
        RECT  2.425 0.940 2.430 2.585 ;
        RECT  1.990 0.940 2.425 1.340 ;
        RECT  1.735 1.975 2.425 2.375 ;
        RECT  1.895 0.880 1.990 1.340 ;
        RECT  1.635 0.635 1.895 1.340 ;
        RECT  1.475 1.975 1.735 2.915 ;
        END
        ANTENNADIFFAREA     1.3988 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.545 0.910 1.805 ;
        RECT  0.125 1.290 0.335 1.805 ;
        END
        ANTENNAGATEAREA     0.2847 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.465 -0.250 3.220 0.250 ;
        RECT  2.205 -0.250 2.465 0.405 ;
        RECT  1.325 -0.250 2.205 0.250 ;
        RECT  1.065 -0.250 1.325 0.965 ;
        RECT  0.000 -0.250 1.065 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.090 3.440 3.220 3.940 ;
        RECT  2.830 3.285 3.090 3.940 ;
        RECT  2.150 3.440 2.830 3.940 ;
        RECT  1.890 3.285 2.150 3.940 ;
        RECT  1.195 3.440 1.890 3.940 ;
        RECT  0.935 3.285 1.195 3.940 ;
        RECT  0.725 3.440 0.935 3.940 ;
        RECT  0.125 3.045 0.725 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.265 1.535 2.245 1.795 ;
        RECT  1.105 1.205 1.265 2.145 ;
        RECT  0.785 1.205 1.105 1.365 ;
        RECT  0.785 1.985 1.105 2.145 ;
        RECT  0.625 0.845 0.785 1.365 ;
        RECT  0.525 1.985 0.785 2.590 ;
        RECT  0.525 0.845 0.625 1.105 ;
    END
END CLKBUFX8

MACRO CLKBUFX6
    CLASS CORE ;
    FOREIGN CLKBUFX6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 1.000 2.635 2.585 ;
        RECT  2.285 1.000 2.545 2.980 ;
        RECT  1.965 1.000 2.285 2.340 ;
        RECT  1.570 1.000 1.965 1.300 ;
        RECT  1.465 2.040 1.965 2.340 ;
        RECT  1.310 0.640 1.570 1.300 ;
        RECT  1.205 2.040 1.465 2.980 ;
        END
        ANTENNADIFFAREA     1.1800 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.545 0.625 1.805 ;
        RECT  0.125 1.545 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2106 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 -0.250 2.760 0.250 ;
        RECT  1.850 -0.250 2.110 0.810 ;
        RECT  1.030 -0.250 1.850 0.250 ;
        RECT  0.770 -0.250 1.030 0.810 ;
        RECT  0.000 -0.250 0.770 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.005 3.440 2.760 3.940 ;
        RECT  1.745 2.555 2.005 3.940 ;
        RECT  0.925 3.440 1.745 3.940 ;
        RECT  0.665 2.555 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.025 1.570 1.740 1.830 ;
        RECT  0.865 1.080 1.025 2.335 ;
        RECT  0.490 1.080 0.865 1.240 ;
        RECT  0.385 2.175 0.865 2.335 ;
        RECT  0.230 0.980 0.490 1.240 ;
        RECT  0.125 2.175 0.385 3.115 ;
    END
END CLKBUFX6

MACRO CLKBUFX4
    CLASS CORE ;
    FOREIGN CLKBUFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 1.090 2.175 2.210 ;
        RECT  1.575 1.090 1.935 1.330 ;
        RECT  1.560 1.970 1.935 2.210 ;
        RECT  1.335 0.850 1.575 1.330 ;
        RECT  1.300 1.970 1.560 3.045 ;
        RECT  1.275 0.850 1.335 1.110 ;
        END
        ANTENNADIFFAREA     0.6574 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.365 1.420 0.625 1.680 ;
        RECT  0.335 1.420 0.365 1.580 ;
        RECT  0.125 1.290 0.335 1.580 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.075 -0.250 2.300 0.250 ;
        RECT  1.815 -0.250 2.075 0.795 ;
        RECT  0.995 -0.250 1.815 0.250 ;
        RECT  0.735 -0.250 0.995 0.745 ;
        RECT  0.000 -0.250 0.735 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 3.440 2.300 3.940 ;
        RECT  1.840 2.555 2.100 3.940 ;
        RECT  1.020 3.440 1.840 3.940 ;
        RECT  0.760 2.215 1.020 3.940 ;
        RECT  0.000 3.440 0.760 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.110 1.510 1.705 1.770 ;
        RECT  1.065 1.510 1.110 2.035 ;
        RECT  0.905 0.950 1.065 2.035 ;
        RECT  0.425 0.950 0.905 1.110 ;
        RECT  0.455 1.875 0.905 2.035 ;
        RECT  0.250 1.875 0.455 2.645 ;
        RECT  0.165 0.850 0.425 1.110 ;
        RECT  0.195 2.045 0.250 2.645 ;
    END
END CLKBUFX4

MACRO CLKBUFX3
    CLASS CORE ;
    FOREIGN CLKBUFX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.690 1.105 1.715 2.175 ;
        RECT  1.535 1.105 1.690 2.220 ;
        RECT  1.505 0.695 1.535 2.220 ;
        RECT  1.275 0.695 1.505 1.295 ;
        RECT  1.295 2.060 1.505 2.220 ;
        RECT  1.035 2.060 1.295 2.660 ;
        END
        ANTENNADIFFAREA     0.5926 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.715 2.110 0.795 2.400 ;
        RECT  0.585 1.265 0.715 2.400 ;
        RECT  0.555 1.265 0.585 2.335 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.995 -0.250 1.840 0.250 ;
        RECT  0.735 -0.250 0.995 0.745 ;
        RECT  0.000 -0.250 0.735 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.695 3.440 1.840 3.940 ;
        RECT  1.435 3.285 1.695 3.940 ;
        RECT  0.895 3.440 1.435 3.940 ;
        RECT  0.635 3.285 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.090 1.550 1.325 1.810 ;
        RECT  0.930 0.925 1.090 1.810 ;
        RECT  0.420 0.925 0.930 1.085 ;
        RECT  0.370 0.825 0.420 1.085 ;
        RECT  0.370 2.835 0.385 3.095 ;
        RECT  0.210 0.825 0.370 3.095 ;
        RECT  0.160 0.825 0.210 1.085 ;
        RECT  0.125 2.835 0.210 3.095 ;
    END
END CLKBUFX3

MACRO CLKBUFX2
    CLASS CORE ;
    FOREIGN CLKBUFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.690 1.105 1.715 2.175 ;
        RECT  1.665 0.920 1.690 2.175 ;
        RECT  1.530 0.920 1.665 2.360 ;
        RECT  1.505 0.820 1.530 2.360 ;
        RECT  1.235 0.820 1.505 1.080 ;
        RECT  1.315 2.200 1.505 2.360 ;
        RECT  1.055 2.200 1.315 2.460 ;
        END
        ANTENNADIFFAREA     0.4130 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.175 0.795 1.680 ;
        RECT  0.455 1.420 0.585 1.680 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 -0.250 1.840 0.250 ;
        RECT  0.695 -0.250 0.955 0.965 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 3.440 1.840 3.940 ;
        RECT  1.455 3.285 1.715 3.940 ;
        RECT  0.825 3.440 1.455 3.940 ;
        RECT  0.565 2.200 0.825 3.940 ;
        RECT  0.545 2.200 0.565 2.460 ;
        RECT  0.000 3.440 0.565 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.225 1.385 1.325 1.645 ;
        RECT  1.065 1.385 1.225 2.020 ;
        RECT  0.285 1.860 1.065 2.020 ;
        RECT  0.275 0.820 0.385 1.080 ;
        RECT  0.285 2.780 0.385 3.040 ;
        RECT  0.275 1.860 0.285 3.040 ;
        RECT  0.115 0.820 0.275 3.040 ;
    END
END CLKBUFX2

MACRO XNOR3X4
    CLASS CORE ;
    FOREIGN XNOR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.165 1.040 11.375 2.395 ;
        RECT  10.915 1.040 11.165 1.250 ;
        RECT  10.915 2.185 11.165 2.395 ;
        RECT  10.845 0.695 10.915 1.250 ;
        RECT  10.865 2.185 10.915 2.995 ;
        RECT  10.605 2.185 10.865 3.125 ;
        RECT  10.635 0.510 10.845 1.250 ;
        RECT  10.575 0.510 10.635 1.110 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.245 1.290 10.455 1.615 ;
        RECT  10.105 1.405 10.245 1.615 ;
        RECT  9.845 1.405 10.105 1.665 ;
        END
        ANTENNAGATEAREA     0.5954 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.235 1.515 6.315 1.990 ;
        RECT  6.130 1.345 6.235 2.300 ;
        RECT  6.075 1.290 6.130 2.300 ;
        RECT  6.015 1.290 6.075 1.505 ;
        RECT  5.755 1.245 6.015 1.505 ;
        END
        ANTENNAGATEAREA     0.9542 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.580 0.425 1.990 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.375 -0.250 11.500 0.250 ;
        RECT  11.115 -0.250 11.375 0.795 ;
        RECT  10.295 -0.250 11.115 0.250 ;
        RECT  10.035 -0.250 10.295 1.105 ;
        RECT  4.305 -0.250 10.035 0.250 ;
        RECT  4.045 -0.250 4.305 0.405 ;
        RECT  3.225 -0.250 4.045 0.250 ;
        RECT  2.965 -0.250 3.225 0.405 ;
        RECT  0.385 -0.250 2.965 0.250 ;
        RECT  0.125 -0.250 0.385 1.285 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.375 3.440 11.500 3.940 ;
        RECT  11.115 2.595 11.375 3.940 ;
        RECT  10.325 3.440 11.115 3.940 ;
        RECT  10.065 2.860 10.325 3.940 ;
        RECT  4.045 3.440 10.065 3.940 ;
        RECT  3.785 3.115 4.045 3.940 ;
        RECT  2.995 3.440 3.785 3.940 ;
        RECT  2.735 2.790 2.995 3.940 ;
        RECT  0.385 3.440 2.735 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.795 1.550 10.895 1.810 ;
        RECT  10.635 1.550 10.795 2.005 ;
        RECT  10.270 1.845 10.635 2.005 ;
        RECT  10.110 1.845 10.270 2.680 ;
        RECT  9.685 2.520 10.110 2.680 ;
        RECT  9.665 0.930 9.785 1.190 ;
        RECT  9.665 2.080 9.785 2.340 ;
        RECT  9.525 2.520 9.685 3.155 ;
        RECT  9.505 0.930 9.665 2.340 ;
        RECT  8.775 2.995 9.525 3.155 ;
        RECT  9.295 1.525 9.505 1.785 ;
        RECT  9.115 0.870 9.275 1.130 ;
        RECT  9.115 2.215 9.225 2.815 ;
        RECT  8.955 0.470 9.115 2.815 ;
        RECT  7.185 0.470 8.955 0.630 ;
        RECT  8.615 0.810 8.775 3.155 ;
        RECT  8.505 0.810 8.615 1.110 ;
        RECT  8.455 2.320 8.615 2.920 ;
        RECT  7.685 0.810 8.505 0.970 ;
        RECT  8.095 1.150 8.225 1.310 ;
        RECT  8.095 2.055 8.205 2.995 ;
        RECT  7.935 1.150 8.095 3.220 ;
        RECT  4.385 3.060 7.935 3.220 ;
        RECT  7.585 2.245 7.695 2.845 ;
        RECT  7.585 0.810 7.685 1.070 ;
        RECT  7.425 0.810 7.585 2.845 ;
        RECT  7.025 0.470 7.185 2.840 ;
        RECT  6.915 0.470 7.025 1.285 ;
        RECT  6.925 2.240 7.025 2.840 ;
        RECT  6.125 0.470 6.915 0.630 ;
        RECT  6.515 0.810 6.675 2.880 ;
        RECT  6.405 0.810 6.515 1.070 ;
        RECT  6.415 2.280 6.515 2.880 ;
        RECT  4.725 2.720 6.415 2.880 ;
        RECT  5.965 0.470 6.125 1.065 ;
        RECT  5.575 0.805 5.965 1.065 ;
        RECT  5.795 2.280 5.895 2.540 ;
        RECT  5.635 1.920 5.795 2.540 ;
        RECT  5.575 1.920 5.635 2.080 ;
        RECT  5.525 0.805 5.575 2.080 ;
        RECT  5.415 0.905 5.525 2.080 ;
        RECT  5.235 2.270 5.385 2.530 ;
        RECT  5.235 0.475 5.245 0.735 ;
        RECT  5.075 0.475 5.235 2.530 ;
        RECT  4.985 0.475 5.075 0.745 ;
        RECT  3.765 0.585 4.985 0.745 ;
        RECT  4.735 0.975 4.895 1.925 ;
        RECT  4.585 0.975 4.735 1.235 ;
        RECT  4.585 1.695 4.735 1.925 ;
        RECT  4.565 2.435 4.725 2.880 ;
        RECT  4.325 1.695 4.585 2.255 ;
        RECT  4.010 2.435 4.565 2.595 ;
        RECT  4.225 2.775 4.385 3.220 ;
        RECT  2.255 1.695 4.325 1.855 ;
        RECT  3.425 2.775 4.225 2.935 ;
        RECT  3.850 2.065 4.010 2.595 ;
        RECT  3.505 2.065 3.850 2.225 ;
        RECT  3.505 0.430 3.765 0.745 ;
        RECT  3.665 0.930 3.765 1.190 ;
        RECT  3.505 0.930 3.665 1.410 ;
        RECT  2.775 0.585 3.505 0.745 ;
        RECT  1.945 1.250 3.505 1.410 ;
        RECT  3.245 2.065 3.505 2.250 ;
        RECT  3.265 2.450 3.425 2.935 ;
        RECT  2.425 2.450 3.265 2.610 ;
        RECT  1.915 2.065 3.245 2.225 ;
        RECT  2.615 0.470 2.775 0.745 ;
        RECT  0.895 0.470 2.615 0.630 ;
        RECT  2.275 0.810 2.435 1.070 ;
        RECT  2.165 2.405 2.425 3.060 ;
        RECT  1.405 0.810 2.275 0.970 ;
        RECT  1.995 1.595 2.255 1.855 ;
        RECT  1.405 2.900 2.165 3.060 ;
        RECT  1.815 1.150 1.945 1.410 ;
        RECT  1.815 2.065 1.915 2.720 ;
        RECT  1.655 1.150 1.815 2.720 ;
        RECT  1.305 0.810 1.405 1.070 ;
        RECT  1.305 2.045 1.405 3.060 ;
        RECT  1.145 0.810 1.305 3.060 ;
        RECT  0.735 0.470 0.895 3.020 ;
        RECT  0.635 0.470 0.735 1.230 ;
        RECT  0.635 2.080 0.735 3.020 ;
    END
END XNOR3X4

MACRO XNOR3X2
    CLASS CORE ;
    FOREIGN XNOR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.995 0.695 8.155 3.045 ;
        RECT  7.895 0.695 7.995 1.295 ;
        RECT  7.895 2.105 7.995 3.045 ;
        END
        ANTENNADIFFAREA     0.7276 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.645 2.110 7.695 2.400 ;
        RECT  7.485 2.110 7.645 2.665 ;
        RECT  7.130 2.505 7.485 2.665 ;
        RECT  6.970 2.505 7.130 2.970 ;
        END
        ANTENNAGATEAREA     0.2964 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.830 2.110 4.935 2.415 ;
        RECT  4.670 1.260 4.830 2.415 ;
        RECT  4.420 1.260 4.670 1.520 ;
        END
        ANTENNAGATEAREA     0.6812 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.560 0.450 1.995 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.570 -0.250 8.280 0.250 ;
        RECT  6.970 -0.250 7.570 0.405 ;
        RECT  2.545 -0.250 6.970 0.250 ;
        RECT  2.385 -0.250 2.545 1.295 ;
        RECT  0.385 -0.250 2.385 0.250 ;
        RECT  0.125 -0.250 0.385 1.075 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.615 3.440 8.280 3.940 ;
        RECT  7.355 2.895 7.615 3.940 ;
        RECT  2.595 3.440 7.355 3.940 ;
        RECT  2.335 3.090 2.595 3.940 ;
        RECT  0.385 3.440 2.335 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.655 1.540 7.810 1.800 ;
        RECT  7.495 0.625 7.655 1.800 ;
        RECT  6.200 0.625 7.495 0.785 ;
        RECT  6.980 2.030 7.210 2.290 ;
        RECT  6.980 1.085 7.180 1.245 ;
        RECT  6.820 1.085 6.980 2.290 ;
        RECT  6.640 2.540 6.760 2.800 ;
        RECT  6.480 0.965 6.640 3.205 ;
        RECT  6.380 0.965 6.480 1.225 ;
        RECT  2.940 3.045 6.480 3.205 ;
        RECT  6.200 2.265 6.300 2.865 ;
        RECT  6.040 0.625 6.200 2.865 ;
        RECT  5.870 0.625 6.040 1.225 ;
        RECT  5.690 2.265 5.790 2.865 ;
        RECT  5.530 1.430 5.690 2.865 ;
        RECT  5.510 1.430 5.530 1.590 ;
        RECT  5.350 0.470 5.510 1.590 ;
        RECT  4.305 0.470 5.350 0.630 ;
        RECT  5.175 1.770 5.335 2.855 ;
        RECT  5.170 1.770 5.175 1.930 ;
        RECT  5.020 2.595 5.175 2.855 ;
        RECT  5.010 0.920 5.170 1.930 ;
        RECT  3.280 2.695 5.020 2.855 ;
        RECT  4.995 0.920 5.010 1.080 ;
        RECT  4.735 0.820 4.995 1.080 ;
        RECT  4.330 1.915 4.490 2.515 ;
        RECT  4.240 1.915 4.330 2.075 ;
        RECT  4.240 0.470 4.305 1.080 ;
        RECT  4.080 0.470 4.240 2.075 ;
        RECT  3.845 2.255 4.025 2.515 ;
        RECT  3.685 0.540 3.845 2.515 ;
        RECT  3.585 0.540 3.685 1.230 ;
        RECT  2.885 0.540 3.585 0.700 ;
        RECT  3.120 2.410 3.280 2.855 ;
        RECT  3.065 0.885 3.225 2.230 ;
        RECT  1.525 2.410 3.120 2.570 ;
        RECT  1.865 2.070 3.065 2.230 ;
        RECT  2.780 2.750 2.940 3.205 ;
        RECT  2.725 0.540 2.885 1.720 ;
        RECT  1.185 2.750 2.780 2.910 ;
        RECT  2.205 1.560 2.725 1.720 ;
        RECT  2.045 0.475 2.205 1.720 ;
        RECT  0.845 0.475 2.045 0.635 ;
        RECT  1.705 0.815 1.865 1.360 ;
        RECT  1.705 1.545 1.865 2.230 ;
        RECT  1.525 1.200 1.705 1.360 ;
        RECT  1.365 1.200 1.525 2.570 ;
        RECT  1.185 0.815 1.405 0.975 ;
        RECT  1.025 0.815 1.185 2.910 ;
        RECT  0.685 0.475 0.845 3.190 ;
    END
END XNOR3X2

MACRO XNOR3X1
    CLASS CORE ;
    FOREIGN XNOR3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 0.980 7.695 2.715 ;
        RECT  7.510 0.980 7.535 1.355 ;
        RECT  7.435 2.105 7.535 2.715 ;
        RECT  7.435 0.980 7.510 1.240 ;
        END
        ANTENNADIFFAREA     0.3672 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 2.520 6.775 3.005 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 1.700 4.600 2.345 ;
        RECT  4.390 1.700 4.440 1.990 ;
        RECT  4.230 1.165 4.390 1.990 ;
        END
        ANTENNAGATEAREA     0.3601 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.505 0.420 2.050 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.610 -0.250 7.820 0.250 ;
        RECT  7.010 -0.250 7.610 0.405 ;
        RECT  1.945 -0.250 7.010 0.250 ;
        RECT  1.685 -0.250 1.945 0.605 ;
        RECT  0.385 -0.250 1.685 0.250 ;
        RECT  0.125 -0.250 0.385 1.220 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.135 3.440 7.820 3.940 ;
        RECT  6.975 2.115 7.135 3.940 ;
        RECT  2.455 3.440 6.975 3.940 ;
        RECT  2.195 3.100 2.455 3.940 ;
        RECT  0.385 3.440 2.195 3.940 ;
        RECT  0.125 2.335 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.200 1.635 7.355 1.895 ;
        RECT  7.195 0.695 7.200 1.895 ;
        RECT  7.040 0.695 7.195 1.795 ;
        RECT  6.760 0.695 7.040 0.855 ;
        RECT  6.600 0.470 6.760 0.855 ;
        RECT  6.485 1.035 6.700 1.315 ;
        RECT  6.485 2.025 6.615 2.285 ;
        RECT  5.630 0.470 6.600 0.630 ;
        RECT  6.440 1.035 6.485 2.285 ;
        RECT  6.325 1.155 6.440 2.285 ;
        RECT  6.140 2.535 6.300 2.795 ;
        RECT  6.140 0.815 6.190 0.975 ;
        RECT  5.980 0.815 6.140 3.220 ;
        RECT  5.930 0.815 5.980 0.975 ;
        RECT  2.855 3.060 5.980 3.220 ;
        RECT  5.630 2.070 5.790 2.880 ;
        RECT  5.470 0.470 5.630 2.230 ;
        RECT  5.120 0.760 5.280 2.880 ;
        RECT  5.070 0.760 5.120 1.025 ;
        RECT  4.910 0.470 5.070 1.025 ;
        RECT  4.780 1.360 4.940 2.880 ;
        RECT  4.150 0.470 4.910 0.630 ;
        RECT  4.730 1.360 4.780 1.520 ;
        RECT  3.370 2.720 4.780 2.880 ;
        RECT  4.570 0.815 4.730 1.520 ;
        RECT  4.400 0.815 4.570 0.975 ;
        RECT  4.060 2.170 4.220 2.535 ;
        RECT  4.050 0.470 4.150 0.735 ;
        RECT  4.050 2.170 4.060 2.330 ;
        RECT  3.890 0.470 4.050 2.330 ;
        RECT  3.550 0.470 3.710 2.535 ;
        RECT  2.285 0.470 3.550 0.630 ;
        RECT  3.210 0.810 3.370 2.880 ;
        RECT  2.625 0.810 3.210 0.970 ;
        RECT  2.870 1.150 3.030 2.575 ;
        RECT  2.815 1.150 2.870 1.410 ;
        RECT  1.525 2.415 2.870 2.575 ;
        RECT  2.695 2.755 2.855 3.220 ;
        RECT  1.185 2.755 2.695 2.915 ;
        RECT  2.465 0.810 2.625 2.235 ;
        RECT  1.865 2.075 2.465 2.235 ;
        RECT  2.125 0.470 2.285 1.725 ;
        RECT  0.895 0.785 2.125 0.945 ;
        RECT  2.080 1.465 2.125 1.725 ;
        RECT  1.865 1.125 1.915 1.285 ;
        RECT  1.705 1.125 1.865 2.235 ;
        RECT  1.655 1.125 1.705 1.285 ;
        RECT  1.365 1.770 1.525 2.575 ;
        RECT  1.305 1.125 1.405 1.285 ;
        RECT  1.185 1.125 1.305 1.560 ;
        RECT  1.145 1.125 1.185 2.915 ;
        RECT  1.025 1.400 1.145 2.915 ;
        RECT  0.785 0.785 0.895 1.220 ;
        RECT  0.785 2.315 0.845 2.915 ;
        RECT  0.735 0.785 0.785 2.915 ;
        RECT  0.625 0.960 0.735 2.915 ;
    END
END XNOR3X1

MACRO XNOR3XL
    CLASS CORE ;
    FOREIGN XNOR3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 0.960 7.695 2.400 ;
        RECT  7.435 0.960 7.535 1.220 ;
        RECT  7.435 2.025 7.535 2.400 ;
        END
        ANTENNADIFFAREA     0.2176 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 2.520 6.775 3.005 ;
        END
        ANTENNAGATEAREA     0.1560 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 1.700 4.600 2.355 ;
        RECT  4.390 1.700 4.440 1.990 ;
        RECT  4.230 1.165 4.390 1.990 ;
        END
        ANTENNAGATEAREA     0.2340 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.505 0.420 2.050 ;
        END
        ANTENNAGATEAREA     0.0780 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.610 -0.250 7.820 0.250 ;
        RECT  7.010 -0.250 7.610 0.405 ;
        RECT  1.975 -0.250 7.010 0.250 ;
        RECT  1.715 -0.250 1.975 0.605 ;
        RECT  0.385 -0.250 1.715 0.250 ;
        RECT  0.125 -0.250 0.385 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.230 3.440 7.820 3.940 ;
        RECT  6.970 2.025 7.230 3.940 ;
        RECT  6.925 2.025 6.970 2.285 ;
        RECT  2.455 3.440 6.970 3.940 ;
        RECT  2.195 3.100 2.455 3.940 ;
        RECT  0.385 3.440 2.195 3.940 ;
        RECT  0.125 2.705 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.200 1.530 7.355 1.795 ;
        RECT  7.040 0.585 7.200 1.795 ;
        RECT  6.760 0.585 7.040 0.745 ;
        RECT  6.600 0.470 6.760 0.745 ;
        RECT  6.485 0.960 6.700 1.315 ;
        RECT  6.485 2.025 6.615 2.285 ;
        RECT  5.630 0.470 6.600 0.630 ;
        RECT  6.440 0.960 6.485 2.285 ;
        RECT  6.325 1.155 6.440 2.285 ;
        RECT  6.140 2.535 6.300 2.795 ;
        RECT  6.090 0.815 6.190 0.975 ;
        RECT  6.090 1.565 6.140 3.220 ;
        RECT  5.980 0.815 6.090 3.220 ;
        RECT  5.930 0.815 5.980 1.725 ;
        RECT  2.855 3.060 5.980 3.220 ;
        RECT  5.630 1.985 5.790 2.795 ;
        RECT  5.470 0.470 5.630 2.145 ;
        RECT  5.120 0.675 5.280 2.795 ;
        RECT  5.070 0.675 5.120 1.025 ;
        RECT  4.910 0.470 5.070 1.025 ;
        RECT  4.780 1.360 4.940 2.875 ;
        RECT  4.150 0.470 4.910 0.630 ;
        RECT  4.730 1.360 4.780 1.520 ;
        RECT  4.560 2.535 4.780 2.875 ;
        RECT  4.570 0.815 4.730 1.520 ;
        RECT  4.400 0.815 4.570 0.975 ;
        RECT  3.370 2.715 4.560 2.875 ;
        RECT  4.060 2.170 4.220 2.535 ;
        RECT  4.050 0.470 4.150 0.735 ;
        RECT  4.050 2.170 4.060 2.330 ;
        RECT  3.890 0.470 4.050 2.330 ;
        RECT  3.550 0.470 3.710 2.535 ;
        RECT  2.315 0.470 3.550 0.630 ;
        RECT  3.210 0.810 3.370 2.875 ;
        RECT  2.655 0.810 3.210 0.970 ;
        RECT  2.870 1.150 3.030 2.575 ;
        RECT  2.835 1.150 2.870 1.410 ;
        RECT  1.525 2.415 2.870 2.575 ;
        RECT  2.695 2.755 2.855 3.220 ;
        RECT  1.185 2.755 2.695 2.915 ;
        RECT  2.495 0.810 2.655 2.235 ;
        RECT  1.865 2.075 2.495 2.235 ;
        RECT  2.155 0.470 2.315 1.725 ;
        RECT  0.895 0.785 2.155 0.945 ;
        RECT  2.080 1.465 2.155 1.725 ;
        RECT  1.845 1.125 1.945 1.285 ;
        RECT  1.845 1.490 1.865 2.235 ;
        RECT  1.705 1.125 1.845 2.235 ;
        RECT  1.685 1.125 1.705 1.650 ;
        RECT  1.365 1.855 1.525 2.575 ;
        RECT  1.305 1.125 1.435 1.285 ;
        RECT  1.185 1.125 1.305 1.675 ;
        RECT  1.145 1.125 1.185 2.915 ;
        RECT  1.025 1.515 1.145 2.915 ;
        RECT  0.785 0.785 0.895 1.295 ;
        RECT  0.785 2.705 0.845 2.965 ;
        RECT  0.735 0.785 0.785 2.965 ;
        RECT  0.625 1.035 0.735 2.965 ;
    END
END XNOR3XL

MACRO XNOR2X4
    CLASS CORE ;
    FOREIGN XNOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.145 0.880 8.155 2.700 ;
        RECT  7.945 0.585 8.145 2.700 ;
        RECT  6.325 0.585 7.945 0.785 ;
        RECT  6.695 2.500 7.945 2.700 ;
        RECT  6.495 2.500 6.695 3.150 ;
        RECT  3.335 2.950 6.495 3.150 ;
        RECT  6.125 0.585 6.325 1.205 ;
        RECT  5.485 1.005 6.125 1.205 ;
        RECT  5.225 0.905 5.485 1.205 ;
        RECT  4.465 1.005 5.225 1.205 ;
        RECT  4.205 0.815 4.465 1.205 ;
        RECT  3.405 0.815 4.205 1.005 ;
        RECT  3.145 0.815 3.405 1.075 ;
        RECT  3.075 2.890 3.335 3.150 ;
        END
        ANTENNADIFFAREA     1.9866 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.595 1.165 1.855 ;
        RECT  0.585 1.595 0.795 1.990 ;
        RECT  0.565 1.595 0.585 1.855 ;
        END
        ANTENNAGATEAREA     0.6318 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 1.595 2.185 1.855 ;
        RECT  1.715 1.595 1.925 1.805 ;
        RECT  1.505 1.290 1.715 1.805 ;
        END
        ANTENNAGATEAREA     0.9308 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.095 -0.250 8.280 0.250 ;
        RECT  7.835 -0.250 8.095 0.405 ;
        RECT  7.115 -0.250 7.835 0.250 ;
        RECT  6.855 -0.250 7.115 0.405 ;
        RECT  1.805 -0.250 6.855 0.250 ;
        RECT  1.545 -0.250 1.805 0.405 ;
        RECT  0.895 -0.250 1.545 0.250 ;
        RECT  0.635 -0.250 0.895 0.945 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.155 3.440 8.280 3.940 ;
        RECT  7.895 2.900 8.155 3.940 ;
        RECT  7.135 3.440 7.895 3.940 ;
        RECT  6.875 2.900 7.135 3.940 ;
        RECT  1.915 3.440 6.875 3.940 ;
        RECT  1.655 2.810 1.915 3.940 ;
        RECT  0.895 3.440 1.655 3.940 ;
        RECT  0.635 2.670 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.505 0.965 7.665 2.320 ;
        RECT  7.405 0.965 7.505 1.225 ;
        RECT  6.365 2.160 7.505 2.320 ;
        RECT  6.665 1.065 7.405 1.225 ;
        RECT  6.935 1.720 7.195 1.980 ;
        RECT  6.180 1.820 6.935 1.980 ;
        RECT  6.505 1.065 6.665 1.545 ;
        RECT  5.835 1.385 6.505 1.545 ;
        RECT  6.020 1.820 6.180 2.765 ;
        RECT  3.845 2.605 6.020 2.765 ;
        RECT  5.785 0.475 5.945 0.825 ;
        RECT  5.675 1.385 5.835 2.425 ;
        RECT  4.975 0.475 5.785 0.635 ;
        RECT  3.955 1.385 5.675 1.545 ;
        RECT  4.865 2.265 5.675 2.425 ;
        RECT  4.435 1.725 5.035 1.985 ;
        RECT  4.715 0.475 4.975 0.825 ;
        RECT  4.605 2.165 4.865 2.425 ;
        RECT  2.145 0.475 4.715 0.635 ;
        RECT  2.530 1.825 4.435 1.985 ;
        RECT  3.695 1.185 3.955 1.545 ;
        RECT  3.585 2.165 3.845 2.765 ;
        RECT  2.960 1.385 3.695 1.545 ;
        RECT  2.825 2.470 3.585 2.630 ;
        RECT  2.800 0.815 2.960 1.545 ;
        RECT  2.565 2.470 2.825 2.830 ;
        RECT  2.635 0.815 2.800 1.075 ;
        RECT  1.405 2.470 2.565 2.630 ;
        RECT  2.370 1.255 2.530 2.270 ;
        RECT  2.355 1.255 2.370 1.415 ;
        RECT  2.165 2.110 2.370 2.270 ;
        RECT  2.095 1.035 2.355 1.415 ;
        RECT  1.985 0.475 2.145 0.835 ;
        RECT  1.405 0.675 1.985 0.835 ;
        RECT  1.295 0.675 1.405 1.075 ;
        RECT  1.145 2.080 1.405 3.020 ;
        RECT  1.135 0.675 1.295 1.285 ;
        RECT  0.385 2.170 1.145 2.330 ;
        RECT  0.385 1.125 1.135 1.285 ;
        RECT  0.285 0.685 0.385 1.285 ;
        RECT  0.285 2.080 0.385 3.020 ;
        RECT  0.125 0.685 0.285 3.020 ;
    END
END XNOR2X4

MACRO XNOR2X2
    CLASS CORE ;
    FOREIGN XNOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.295 0.845 5.395 2.755 ;
        RECT  5.135 0.585 5.295 2.755 ;
        RECT  4.375 0.585 5.135 0.745 ;
        RECT  4.215 0.585 4.375 2.755 ;
        RECT  4.115 0.585 4.215 1.105 ;
        RECT  4.115 2.155 4.215 2.755 ;
        RECT  3.355 0.585 4.115 0.745 ;
        RECT  3.195 0.585 3.355 2.415 ;
        RECT  3.095 0.815 3.195 1.075 ;
        RECT  3.095 2.155 3.195 2.415 ;
        END
        ANTENNADIFFAREA     1.3780 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.370 0.990 1.630 ;
        RECT  0.585 1.290 0.795 1.630 ;
        RECT  0.390 1.370 0.585 1.630 ;
        END
        ANTENNAGATEAREA     0.3380 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.630 2.500 2.025 ;
        END
        ANTENNAGATEAREA     0.4693 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 -0.250 5.520 0.250 ;
        RECT  2.110 -0.250 2.370 0.405 ;
        RECT  1.335 -0.250 2.110 0.250 ;
        RECT  1.075 -0.250 1.335 0.405 ;
        RECT  0.385 -0.250 1.075 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.255 3.440 5.520 3.940 ;
        RECT  1.995 3.285 2.255 3.940 ;
        RECT  1.240 3.440 1.995 3.940 ;
        RECT  0.980 3.285 1.240 3.940 ;
        RECT  0.385 3.440 0.980 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.785 0.925 4.885 1.185 ;
        RECT  4.785 2.175 4.885 2.775 ;
        RECT  4.625 0.925 4.785 3.100 ;
        RECT  1.340 2.940 4.625 3.100 ;
        RECT  3.705 0.925 3.865 2.755 ;
        RECT  3.605 0.925 3.705 1.185 ;
        RECT  3.605 2.155 3.705 2.755 ;
        RECT  1.785 2.595 3.605 2.755 ;
        RECT  2.915 1.685 3.015 1.945 ;
        RECT  2.755 0.945 2.915 2.400 ;
        RECT  2.585 0.945 2.755 1.205 ;
        RECT  2.555 2.240 2.755 2.400 ;
        RECT  1.785 0.935 1.820 1.195 ;
        RECT  1.625 0.935 1.785 2.755 ;
        RECT  1.560 0.935 1.625 1.195 ;
        RECT  1.520 2.115 1.625 2.755 ;
        RECT  1.340 1.410 1.445 1.685 ;
        RECT  1.330 1.410 1.340 3.100 ;
        RECT  1.180 0.925 1.330 3.100 ;
        RECT  1.170 0.925 1.180 2.630 ;
        RECT  0.820 0.925 1.170 1.085 ;
        RECT  0.820 2.395 1.170 2.630 ;
        RECT  0.560 0.825 0.820 1.085 ;
        RECT  0.560 2.130 0.820 2.830 ;
    END
END XNOR2X2

MACRO XNOR2X1
    CLASS CORE ;
    FOREIGN XNOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.075 1.515 2.175 1.990 ;
        RECT  2.060 1.515 2.075 2.420 ;
        RECT  1.900 0.895 2.060 2.420 ;
        RECT  1.800 0.895 1.900 1.155 ;
        RECT  1.815 2.160 1.900 2.420 ;
        END
        ANTENNADIFFAREA     0.5036 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.970 1.290 1.255 1.850 ;
        END
        ANTENNAGATEAREA     0.1690 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.380 1.765 0.430 2.025 ;
        RECT  0.100 1.700 0.380 2.205 ;
        END
        ANTENNAGATEAREA     0.2340 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 -0.250 3.220 0.250 ;
        RECT  2.820 -0.250 3.080 0.990 ;
        RECT  1.035 -0.250 2.820 0.250 ;
        RECT  0.775 -0.250 1.035 0.990 ;
        RECT  0.000 -0.250 0.775 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.045 3.440 3.220 3.940 ;
        RECT  2.885 2.085 3.045 3.940 ;
        RECT  0.935 3.440 2.885 3.940 ;
        RECT  0.675 2.950 0.935 3.940 ;
        RECT  0.000 3.440 0.675 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.520 2.625 2.680 3.170 ;
        RECT  2.570 2.160 2.585 2.420 ;
        RECT  2.410 0.895 2.570 2.420 ;
        RECT  1.630 2.625 2.520 2.785 ;
        RECT  2.310 0.895 2.410 1.155 ;
        RECT  2.325 2.160 2.410 2.420 ;
        RECT  1.985 2.975 2.245 3.185 ;
        RECT  1.290 2.975 1.985 3.135 ;
        RECT  1.595 2.210 1.630 2.785 ;
        RECT  1.470 0.800 1.595 2.785 ;
        RECT  1.435 0.800 1.470 2.420 ;
        RECT  1.290 0.800 1.435 1.060 ;
        RECT  1.305 2.160 1.435 2.420 ;
        RECT  1.130 2.605 1.290 3.135 ;
        RECT  0.770 2.605 1.130 2.765 ;
        RECT  0.610 1.330 0.770 2.765 ;
        RECT  0.445 1.330 0.610 1.490 ;
        RECT  0.125 2.425 0.610 2.685 ;
        RECT  0.285 0.950 0.445 1.490 ;
        RECT  0.185 0.950 0.285 1.210 ;
    END
END XNOR2X1

MACRO XNOR2XL
    CLASS CORE ;
    FOREIGN XNOR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.030 2.270 2.745 ;
        RECT  2.110 1.030 2.175 3.220 ;
        RECT  2.095 1.030 2.110 1.190 ;
        RECT  2.015 2.585 2.110 3.220 ;
        RECT  1.835 0.930 2.095 1.190 ;
        RECT  1.835 2.585 2.015 2.745 ;
        RECT  1.965 2.930 2.015 3.220 ;
        END
        ANTENNADIFFAREA     0.2377 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.465 1.090 1.725 ;
        RECT  0.585 1.290 0.795 1.725 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.790 0.500 3.140 ;
        RECT  0.125 2.790 0.335 3.220 ;
        RECT  0.120 2.790 0.125 3.140 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.220 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.955 -0.250 2.835 0.250 ;
        RECT  0.695 -0.250 0.955 1.110 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.220 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.955 3.440 2.835 3.940 ;
        RECT  0.695 2.335 0.955 3.940 ;
        RECT  0.000 3.440 0.695 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.805 0.590 2.965 1.735 ;
        RECT  1.580 0.590 2.805 0.750 ;
        RECT  2.455 0.930 2.615 2.705 ;
        RECT  1.770 1.400 1.930 2.405 ;
        RECT  1.580 1.400 1.770 1.560 ;
        RECT  1.525 2.245 1.770 2.405 ;
        RECT  1.430 1.785 1.590 2.065 ;
        RECT  1.420 0.590 1.580 1.560 ;
        RECT  1.265 2.245 1.525 2.595 ;
        RECT  0.385 1.905 1.430 2.065 ;
        RECT  1.265 0.930 1.420 1.190 ;
        RECT  0.285 0.915 0.385 1.175 ;
        RECT  0.285 1.905 0.385 2.485 ;
        RECT  0.125 0.915 0.285 2.485 ;
    END
END XNOR2XL

MACRO XOR3X4
    CLASS CORE ;
    FOREIGN XOR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.165 1.040 11.375 2.395 ;
        RECT  10.915 1.040 11.165 1.250 ;
        RECT  10.915 2.185 11.165 2.395 ;
        RECT  10.845 0.695 10.915 1.250 ;
        RECT  10.865 2.185 10.915 2.995 ;
        RECT  10.605 2.185 10.865 3.125 ;
        RECT  10.635 0.510 10.845 1.250 ;
        RECT  10.575 0.510 10.635 1.110 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.245 1.290 10.455 1.615 ;
        RECT  10.105 1.405 10.245 1.615 ;
        RECT  9.845 1.405 10.105 1.665 ;
        END
        ANTENNAGATEAREA     0.5993 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.235 1.515 6.315 1.990 ;
        RECT  6.130 1.345 6.235 2.300 ;
        RECT  6.075 1.290 6.130 2.300 ;
        RECT  6.015 1.290 6.075 1.505 ;
        RECT  5.755 1.245 6.015 1.505 ;
        END
        ANTENNAGATEAREA     0.9542 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.580 0.425 1.990 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.375 -0.250 11.500 0.250 ;
        RECT  11.115 -0.250 11.375 0.795 ;
        RECT  10.295 -0.250 11.115 0.250 ;
        RECT  10.035 -0.250 10.295 1.025 ;
        RECT  4.305 -0.250 10.035 0.250 ;
        RECT  4.045 -0.250 4.305 0.405 ;
        RECT  3.225 -0.250 4.045 0.250 ;
        RECT  2.965 -0.250 3.225 0.405 ;
        RECT  0.385 -0.250 2.965 0.250 ;
        RECT  0.125 -0.250 0.385 1.285 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.375 3.440 11.500 3.940 ;
        RECT  11.115 2.595 11.375 3.940 ;
        RECT  10.325 3.440 11.115 3.940 ;
        RECT  10.065 2.860 10.325 3.940 ;
        RECT  4.045 3.440 10.065 3.940 ;
        RECT  3.785 3.115 4.045 3.940 ;
        RECT  2.995 3.440 3.785 3.940 ;
        RECT  2.735 2.790 2.995 3.940 ;
        RECT  0.385 3.440 2.735 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.795 1.550 10.895 1.810 ;
        RECT  10.635 1.550 10.795 2.005 ;
        RECT  10.270 1.845 10.635 2.005 ;
        RECT  10.110 1.845 10.270 2.680 ;
        RECT  9.685 2.520 10.110 2.680 ;
        RECT  9.635 2.080 9.785 2.340 ;
        RECT  9.635 0.930 9.755 1.190 ;
        RECT  9.525 2.520 9.685 3.060 ;
        RECT  9.475 0.930 9.635 2.340 ;
        RECT  8.715 2.900 9.525 3.060 ;
        RECT  9.295 1.555 9.475 1.815 ;
        RECT  9.115 2.110 9.225 2.710 ;
        RECT  9.115 0.470 9.215 0.785 ;
        RECT  8.955 0.470 9.115 2.710 ;
        RECT  7.185 0.470 8.955 0.630 ;
        RECT  8.555 0.810 8.715 3.060 ;
        RECT  8.445 0.810 8.555 1.110 ;
        RECT  8.455 2.320 8.555 3.060 ;
        RECT  7.685 0.810 8.445 0.970 ;
        RECT  8.095 2.245 8.205 3.220 ;
        RECT  8.095 1.150 8.195 1.310 ;
        RECT  7.935 1.150 8.095 3.220 ;
        RECT  4.385 3.060 7.935 3.220 ;
        RECT  7.585 2.245 7.695 2.845 ;
        RECT  7.585 0.810 7.685 1.070 ;
        RECT  7.425 0.810 7.585 2.845 ;
        RECT  7.025 0.470 7.185 2.840 ;
        RECT  6.915 0.470 7.025 1.295 ;
        RECT  6.925 2.240 7.025 2.840 ;
        RECT  6.125 0.470 6.915 0.630 ;
        RECT  6.515 0.810 6.675 2.880 ;
        RECT  6.405 0.810 6.515 1.070 ;
        RECT  6.415 2.280 6.515 2.880 ;
        RECT  4.725 2.720 6.415 2.880 ;
        RECT  5.965 0.470 6.125 1.065 ;
        RECT  5.575 0.805 5.965 1.065 ;
        RECT  5.795 2.280 5.895 2.540 ;
        RECT  5.635 1.920 5.795 2.540 ;
        RECT  5.575 1.920 5.635 2.080 ;
        RECT  5.525 0.805 5.575 2.080 ;
        RECT  5.415 0.905 5.525 2.080 ;
        RECT  5.235 2.270 5.385 2.530 ;
        RECT  5.235 0.475 5.245 0.735 ;
        RECT  5.075 0.475 5.235 2.530 ;
        RECT  4.985 0.475 5.075 0.745 ;
        RECT  3.765 0.585 4.985 0.745 ;
        RECT  4.735 0.975 4.895 1.925 ;
        RECT  4.585 0.975 4.735 1.235 ;
        RECT  4.585 1.695 4.735 1.925 ;
        RECT  4.565 2.435 4.725 2.880 ;
        RECT  4.325 1.695 4.585 2.255 ;
        RECT  4.010 2.435 4.565 2.595 ;
        RECT  4.225 2.775 4.385 3.220 ;
        RECT  2.255 1.695 4.325 1.855 ;
        RECT  3.425 2.775 4.225 2.935 ;
        RECT  3.850 2.065 4.010 2.595 ;
        RECT  3.505 2.065 3.850 2.225 ;
        RECT  3.505 0.430 3.765 0.745 ;
        RECT  3.665 0.930 3.765 1.190 ;
        RECT  3.505 0.930 3.665 1.410 ;
        RECT  2.775 0.585 3.505 0.745 ;
        RECT  1.945 1.250 3.505 1.410 ;
        RECT  3.245 2.065 3.505 2.250 ;
        RECT  3.265 2.450 3.425 2.935 ;
        RECT  2.425 2.450 3.265 2.610 ;
        RECT  1.915 2.065 3.245 2.225 ;
        RECT  2.615 0.470 2.775 0.745 ;
        RECT  0.895 0.470 2.615 0.630 ;
        RECT  2.275 0.810 2.435 1.070 ;
        RECT  2.165 2.405 2.425 3.060 ;
        RECT  1.405 0.810 2.275 0.970 ;
        RECT  1.995 1.595 2.255 1.855 ;
        RECT  1.405 2.900 2.165 3.060 ;
        RECT  1.815 1.150 1.945 1.410 ;
        RECT  1.815 2.065 1.915 2.720 ;
        RECT  1.655 1.150 1.815 2.720 ;
        RECT  1.305 0.810 1.405 1.070 ;
        RECT  1.305 2.045 1.405 3.060 ;
        RECT  1.145 0.810 1.305 3.060 ;
        RECT  0.735 0.470 0.895 3.020 ;
        RECT  0.635 0.470 0.735 1.230 ;
        RECT  0.635 2.080 0.735 3.020 ;
    END
END XOR3X4

MACRO XOR3X2
    CLASS CORE ;
    FOREIGN XOR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.995 0.695 8.155 3.045 ;
        RECT  7.895 0.695 7.995 1.295 ;
        RECT  7.895 2.105 7.995 3.045 ;
        END
        ANTENNADIFFAREA     0.7276 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.645 2.110 7.695 2.400 ;
        RECT  7.485 2.110 7.645 2.665 ;
        RECT  7.145 2.505 7.485 2.665 ;
        RECT  6.985 2.505 7.145 2.885 ;
        END
        ANTENNAGATEAREA     0.2990 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.830 2.110 4.935 2.420 ;
        RECT  4.670 1.260 4.830 2.420 ;
        RECT  4.420 1.260 4.670 1.520 ;
        END
        ANTENNAGATEAREA     0.6812 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.560 0.450 1.995 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.570 -0.250 8.280 0.250 ;
        RECT  6.970 -0.250 7.570 0.405 ;
        RECT  2.545 -0.250 6.970 0.250 ;
        RECT  2.385 -0.250 2.545 1.295 ;
        RECT  0.385 -0.250 2.385 0.250 ;
        RECT  0.125 -0.250 0.385 1.075 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.615 3.440 8.280 3.940 ;
        RECT  7.355 2.895 7.615 3.940 ;
        RECT  2.595 3.440 7.355 3.940 ;
        RECT  2.335 3.090 2.595 3.940 ;
        RECT  0.385 3.440 2.335 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.655 1.540 7.810 1.800 ;
        RECT  7.495 0.695 7.655 1.800 ;
        RECT  6.200 0.695 7.495 0.855 ;
        RECT  6.980 2.030 7.210 2.290 ;
        RECT  6.980 1.085 7.180 1.245 ;
        RECT  6.820 1.085 6.980 2.290 ;
        RECT  6.640 2.540 6.760 2.800 ;
        RECT  6.480 1.035 6.640 3.205 ;
        RECT  6.380 1.035 6.480 1.295 ;
        RECT  2.940 3.045 6.480 3.205 ;
        RECT  6.200 2.265 6.300 2.865 ;
        RECT  6.040 0.695 6.200 2.865 ;
        RECT  5.870 0.695 6.040 1.295 ;
        RECT  5.690 2.265 5.790 2.865 ;
        RECT  5.570 1.430 5.690 2.865 ;
        RECT  5.530 0.470 5.570 2.865 ;
        RECT  5.410 0.470 5.530 1.590 ;
        RECT  4.305 0.470 5.410 0.630 ;
        RECT  5.220 1.770 5.335 2.860 ;
        RECT  5.175 0.920 5.220 2.860 ;
        RECT  5.060 0.920 5.175 1.930 ;
        RECT  5.020 2.600 5.175 2.860 ;
        RECT  4.995 0.920 5.060 1.080 ;
        RECT  3.280 2.700 5.020 2.860 ;
        RECT  4.735 0.820 4.995 1.080 ;
        RECT  4.330 1.915 4.490 2.515 ;
        RECT  4.240 1.915 4.330 2.075 ;
        RECT  4.240 0.470 4.305 1.080 ;
        RECT  4.080 0.470 4.240 2.075 ;
        RECT  3.845 2.255 4.025 2.515 ;
        RECT  3.685 0.540 3.845 2.515 ;
        RECT  3.585 0.540 3.685 1.230 ;
        RECT  2.885 0.540 3.585 0.700 ;
        RECT  3.120 2.410 3.280 2.860 ;
        RECT  3.065 0.885 3.225 2.230 ;
        RECT  1.525 2.410 3.120 2.570 ;
        RECT  1.865 2.070 3.065 2.230 ;
        RECT  2.780 2.750 2.940 3.205 ;
        RECT  2.725 0.540 2.885 1.720 ;
        RECT  1.185 2.750 2.780 2.910 ;
        RECT  2.205 1.560 2.725 1.720 ;
        RECT  2.045 0.475 2.205 1.720 ;
        RECT  0.845 0.475 2.045 0.635 ;
        RECT  1.705 0.815 1.865 1.360 ;
        RECT  1.705 1.545 1.865 2.230 ;
        RECT  1.525 1.200 1.705 1.360 ;
        RECT  1.365 1.200 1.525 2.570 ;
        RECT  1.185 0.815 1.405 0.975 ;
        RECT  1.025 0.815 1.185 2.910 ;
        RECT  0.685 0.475 0.845 3.190 ;
    END
END XOR3X2

MACRO XOR3X1
    CLASS CORE ;
    FOREIGN XOR3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 0.980 7.695 2.715 ;
        RECT  7.510 0.980 7.535 1.355 ;
        RECT  7.435 2.105 7.535 2.715 ;
        RECT  7.435 0.980 7.510 1.240 ;
        END
        ANTENNADIFFAREA     0.3672 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 2.520 6.775 3.005 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 1.700 4.600 2.345 ;
        RECT  4.390 1.700 4.440 1.990 ;
        RECT  4.230 1.165 4.390 1.990 ;
        END
        ANTENNAGATEAREA     0.3601 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.505 0.420 2.050 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.610 -0.250 7.820 0.250 ;
        RECT  7.010 -0.250 7.610 0.405 ;
        RECT  1.945 -0.250 7.010 0.250 ;
        RECT  1.685 -0.250 1.945 0.605 ;
        RECT  0.385 -0.250 1.685 0.250 ;
        RECT  0.125 -0.250 0.385 1.220 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.135 3.440 7.820 3.940 ;
        RECT  6.975 2.115 7.135 3.940 ;
        RECT  2.455 3.440 6.975 3.940 ;
        RECT  2.195 3.100 2.455 3.940 ;
        RECT  0.385 3.440 2.195 3.940 ;
        RECT  0.125 2.335 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.200 1.635 7.355 1.895 ;
        RECT  7.195 0.695 7.200 1.895 ;
        RECT  7.040 0.695 7.195 1.795 ;
        RECT  6.760 0.695 7.040 0.855 ;
        RECT  6.600 0.470 6.760 0.855 ;
        RECT  6.485 1.035 6.700 1.315 ;
        RECT  6.485 2.025 6.615 2.285 ;
        RECT  5.630 0.470 6.600 0.630 ;
        RECT  6.440 1.035 6.485 2.285 ;
        RECT  6.325 1.155 6.440 2.285 ;
        RECT  6.140 2.535 6.300 2.795 ;
        RECT  6.140 0.815 6.190 0.975 ;
        RECT  5.980 0.815 6.140 3.220 ;
        RECT  5.930 0.815 5.980 0.975 ;
        RECT  2.855 3.060 5.980 3.220 ;
        RECT  5.630 2.070 5.790 2.880 ;
        RECT  5.470 0.470 5.630 2.230 ;
        RECT  5.120 0.760 5.280 2.880 ;
        RECT  5.070 0.760 5.120 1.025 ;
        RECT  4.910 0.470 5.070 1.025 ;
        RECT  4.780 1.360 4.940 2.880 ;
        RECT  4.150 0.470 4.910 0.630 ;
        RECT  4.730 1.360 4.780 1.520 ;
        RECT  3.370 2.720 4.780 2.880 ;
        RECT  4.570 0.815 4.730 1.520 ;
        RECT  4.400 0.815 4.570 0.975 ;
        RECT  4.060 2.170 4.220 2.535 ;
        RECT  4.050 0.470 4.150 0.735 ;
        RECT  4.050 2.170 4.060 2.330 ;
        RECT  3.890 0.470 4.050 2.330 ;
        RECT  3.550 0.470 3.710 2.535 ;
        RECT  2.285 0.470 3.550 0.630 ;
        RECT  3.210 0.810 3.370 2.880 ;
        RECT  2.625 0.810 3.210 0.970 ;
        RECT  2.870 1.150 3.030 2.575 ;
        RECT  2.815 1.150 2.870 1.410 ;
        RECT  1.525 2.415 2.870 2.575 ;
        RECT  2.695 2.755 2.855 3.220 ;
        RECT  1.185 2.755 2.695 2.915 ;
        RECT  2.465 0.810 2.625 2.235 ;
        RECT  1.865 2.075 2.465 2.235 ;
        RECT  2.125 0.470 2.285 1.725 ;
        RECT  0.895 0.785 2.125 0.945 ;
        RECT  2.080 1.465 2.125 1.725 ;
        RECT  1.865 1.125 1.915 1.285 ;
        RECT  1.705 1.125 1.865 2.235 ;
        RECT  1.655 1.125 1.705 1.285 ;
        RECT  1.365 1.770 1.525 2.575 ;
        RECT  1.305 1.125 1.405 1.285 ;
        RECT  1.185 1.125 1.305 1.560 ;
        RECT  1.145 1.125 1.185 2.915 ;
        RECT  1.025 1.400 1.145 2.915 ;
        RECT  0.785 0.785 0.895 1.220 ;
        RECT  0.785 2.315 0.845 2.915 ;
        RECT  0.735 0.785 0.785 2.915 ;
        RECT  0.625 0.960 0.735 2.915 ;
    END
END XOR3X1

MACRO XOR3XL
    CLASS CORE ;
    FOREIGN XOR3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 0.960 7.695 2.400 ;
        RECT  7.435 0.960 7.535 1.220 ;
        RECT  7.435 2.025 7.535 2.400 ;
        END
        ANTENNADIFFAREA     0.2176 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 2.520 6.775 3.005 ;
        END
        ANTENNAGATEAREA     0.1560 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 1.700 4.600 2.355 ;
        RECT  4.390 1.700 4.440 1.990 ;
        RECT  4.230 1.165 4.390 1.990 ;
        END
        ANTENNAGATEAREA     0.2340 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.505 0.420 2.050 ;
        END
        ANTENNAGATEAREA     0.0780 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.610 -0.250 7.820 0.250 ;
        RECT  7.010 -0.250 7.610 0.405 ;
        RECT  1.975 -0.250 7.010 0.250 ;
        RECT  1.715 -0.250 1.975 0.605 ;
        RECT  0.385 -0.250 1.715 0.250 ;
        RECT  0.125 -0.250 0.385 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.230 3.440 7.820 3.940 ;
        RECT  6.970 2.025 7.230 3.940 ;
        RECT  6.925 2.025 6.970 2.285 ;
        RECT  2.455 3.440 6.970 3.940 ;
        RECT  2.195 3.100 2.455 3.940 ;
        RECT  0.385 3.440 2.195 3.940 ;
        RECT  0.125 2.705 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.200 1.530 7.355 1.795 ;
        RECT  7.040 0.585 7.200 1.795 ;
        RECT  6.760 0.585 7.040 0.745 ;
        RECT  6.600 0.470 6.760 0.745 ;
        RECT  6.485 0.960 6.700 1.315 ;
        RECT  6.485 2.025 6.615 2.285 ;
        RECT  5.630 0.470 6.600 0.630 ;
        RECT  6.440 0.960 6.485 2.285 ;
        RECT  6.325 1.155 6.440 2.285 ;
        RECT  6.140 2.535 6.300 2.795 ;
        RECT  6.090 0.815 6.190 0.975 ;
        RECT  6.090 1.440 6.140 3.220 ;
        RECT  5.980 0.815 6.090 3.220 ;
        RECT  5.930 0.815 5.980 1.600 ;
        RECT  2.855 3.060 5.980 3.220 ;
        RECT  5.630 1.985 5.790 2.795 ;
        RECT  5.470 0.470 5.630 2.145 ;
        RECT  5.120 0.675 5.280 2.795 ;
        RECT  5.070 0.675 5.120 1.025 ;
        RECT  4.910 0.470 5.070 1.025 ;
        RECT  4.780 1.360 4.940 2.875 ;
        RECT  4.150 0.470 4.910 0.630 ;
        RECT  4.730 1.360 4.780 1.520 ;
        RECT  4.560 2.535 4.780 2.875 ;
        RECT  4.570 0.815 4.730 1.520 ;
        RECT  4.400 0.815 4.570 0.975 ;
        RECT  3.370 2.715 4.560 2.875 ;
        RECT  4.060 2.170 4.220 2.535 ;
        RECT  4.050 0.470 4.150 0.735 ;
        RECT  4.050 2.170 4.060 2.330 ;
        RECT  3.890 0.470 4.050 2.330 ;
        RECT  3.550 0.470 3.710 2.535 ;
        RECT  2.315 0.470 3.550 0.630 ;
        RECT  3.210 0.810 3.370 2.875 ;
        RECT  2.655 0.810 3.210 0.970 ;
        RECT  2.870 1.150 3.030 2.575 ;
        RECT  2.835 1.150 2.870 1.410 ;
        RECT  1.525 2.415 2.870 2.575 ;
        RECT  2.695 2.755 2.855 3.220 ;
        RECT  1.185 2.755 2.695 2.915 ;
        RECT  2.495 0.810 2.655 2.235 ;
        RECT  1.865 2.075 2.495 2.235 ;
        RECT  2.155 0.470 2.315 1.725 ;
        RECT  0.895 0.785 2.155 0.945 ;
        RECT  2.080 1.465 2.155 1.725 ;
        RECT  1.845 1.125 1.945 1.285 ;
        RECT  1.845 1.485 1.865 2.235 ;
        RECT  1.705 1.125 1.845 2.235 ;
        RECT  1.685 1.125 1.705 1.645 ;
        RECT  1.365 1.855 1.525 2.575 ;
        RECT  1.305 1.125 1.435 1.285 ;
        RECT  1.185 1.125 1.305 1.675 ;
        RECT  1.145 1.125 1.185 2.915 ;
        RECT  1.025 1.515 1.145 2.915 ;
        RECT  0.785 0.785 0.895 1.295 ;
        RECT  0.785 2.705 0.845 2.965 ;
        RECT  0.735 0.785 0.785 2.965 ;
        RECT  0.625 1.035 0.735 2.965 ;
    END
END XOR3XL

MACRO XOR2X4
    CLASS CORE ;
    FOREIGN XOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.725 0.540 5.985 1.140 ;
        RECT  4.965 0.540 5.725 0.700 ;
        RECT  5.440 2.185 5.700 2.475 ;
        RECT  4.750 2.185 5.440 2.425 ;
        RECT  4.705 0.540 4.965 1.220 ;
        RECT  4.680 2.110 4.750 2.425 ;
        RECT  4.560 0.980 4.705 1.220 ;
        RECT  4.560 2.110 4.680 2.475 ;
        RECT  4.420 0.980 4.560 2.475 ;
        RECT  4.265 0.980 4.420 2.425 ;
        RECT  3.945 0.980 4.265 1.220 ;
        RECT  3.660 2.185 4.265 2.425 ;
        RECT  3.685 0.930 3.945 1.220 ;
        RECT  3.400 2.185 3.660 2.475 ;
        END
        ANTENNADIFFAREA     1.9722 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.685 0.960 1.845 ;
        RECT  0.585 1.685 0.795 1.990 ;
        RECT  0.360 1.685 0.585 1.845 ;
        END
        ANTENNAGATEAREA     0.6760 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.245 1.635 2.505 1.895 ;
        RECT  2.175 1.700 2.245 1.895 ;
        RECT  1.965 1.700 2.175 1.990 ;
        END
        ANTENNAGATEAREA     0.9334 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.110 -0.250 8.280 0.250 ;
        RECT  7.850 -0.250 8.110 1.140 ;
        RECT  7.045 -0.250 7.850 0.250 ;
        RECT  6.785 -0.250 7.045 0.830 ;
        RECT  2.355 -0.250 6.785 0.250 ;
        RECT  2.095 -0.250 2.355 0.405 ;
        RECT  1.295 -0.250 2.095 0.250 ;
        RECT  1.035 -0.250 1.295 1.070 ;
        RECT  0.385 -0.250 1.035 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.150 3.440 8.280 3.940 ;
        RECT  7.890 3.285 8.150 3.940 ;
        RECT  7.350 3.440 7.890 3.940 ;
        RECT  7.090 3.285 7.350 3.940 ;
        RECT  2.200 3.440 7.090 3.940 ;
        RECT  1.940 3.285 2.200 3.940 ;
        RECT  1.295 3.440 1.940 3.940 ;
        RECT  1.035 2.570 1.295 3.940 ;
        RECT  0.385 3.440 1.035 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.600 1.975 7.750 2.915 ;
        RECT  7.490 0.590 7.600 2.915 ;
        RECT  7.440 0.590 7.490 2.295 ;
        RECT  7.340 0.590 7.440 1.250 ;
        RECT  6.750 2.135 7.440 2.295 ;
        RECT  6.495 1.090 7.340 1.250 ;
        RECT  6.745 1.565 7.185 1.825 ;
        RECT  6.590 2.135 6.750 2.855 ;
        RECT  6.585 1.565 6.745 1.900 ;
        RECT  6.405 1.740 6.585 1.900 ;
        RECT  6.395 0.590 6.495 1.250 ;
        RECT  6.245 1.740 6.405 3.165 ;
        RECT  6.235 0.590 6.395 1.500 ;
        RECT  5.140 3.005 6.245 3.165 ;
        RECT  6.065 1.340 6.235 1.500 ;
        RECT  5.905 1.340 6.065 2.825 ;
        RECT  5.475 1.340 5.905 1.500 ;
        RECT  4.170 2.665 5.905 2.825 ;
        RECT  5.215 0.925 5.475 1.500 ;
        RECT  4.930 3.005 5.140 3.220 ;
        RECT  2.565 3.060 4.930 3.220 ;
        RECT  4.195 0.540 4.455 0.800 ;
        RECT  3.435 0.540 4.195 0.700 ;
        RECT  3.910 2.615 4.170 2.875 ;
        RECT  2.890 2.715 3.910 2.875 ;
        RECT  3.175 0.540 3.435 1.140 ;
        RECT  2.905 1.500 3.295 1.760 ;
        RECT  1.805 0.625 3.175 0.785 ;
        RECT  2.745 0.985 2.905 2.415 ;
        RECT  2.645 0.985 2.745 1.245 ;
        RECT  2.490 2.155 2.745 2.415 ;
        RECT  2.405 2.670 2.565 3.220 ;
        RECT  1.805 2.670 2.405 2.830 ;
        RECT  1.705 0.625 1.805 1.195 ;
        RECT  1.705 2.180 1.805 2.830 ;
        RECT  1.645 0.625 1.705 2.830 ;
        RECT  1.545 0.935 1.645 2.830 ;
        RECT  0.785 1.280 1.545 1.440 ;
        RECT  0.785 2.210 1.545 2.370 ;
        RECT  0.625 0.890 0.785 1.440 ;
        RECT  0.525 2.210 0.785 2.810 ;
        RECT  0.525 0.890 0.625 1.150 ;
    END
END XOR2X4

MACRO XOR2X2
    CLASS CORE ;
    FOREIGN XOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.295 0.845 5.395 2.755 ;
        RECT  5.135 0.585 5.295 2.755 ;
        RECT  4.375 0.585 5.135 0.745 ;
        RECT  4.215 0.585 4.375 2.755 ;
        RECT  4.115 0.585 4.215 1.105 ;
        RECT  4.115 2.155 4.215 2.755 ;
        RECT  3.355 0.585 4.115 0.745 ;
        RECT  3.195 0.585 3.355 2.415 ;
        RECT  3.095 0.815 3.195 1.075 ;
        RECT  3.095 2.155 3.195 2.415 ;
        END
        ANTENNADIFFAREA     1.3780 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.370 0.990 1.630 ;
        RECT  0.585 1.290 0.795 1.630 ;
        RECT  0.390 1.370 0.585 1.630 ;
        END
        ANTENNAGATEAREA     0.3380 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.630 2.500 2.025 ;
        END
        ANTENNAGATEAREA     0.4693 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 -0.250 5.520 0.250 ;
        RECT  2.110 -0.250 2.370 0.405 ;
        RECT  1.360 -0.250 2.110 0.250 ;
        RECT  1.100 -0.250 1.360 0.405 ;
        RECT  0.420 -0.250 1.100 0.250 ;
        RECT  0.160 -0.250 0.420 0.405 ;
        RECT  0.000 -0.250 0.160 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.255 3.440 5.520 3.940 ;
        RECT  1.995 3.285 2.255 3.940 ;
        RECT  1.240 3.440 1.995 3.940 ;
        RECT  0.980 3.285 1.240 3.940 ;
        RECT  0.420 3.440 0.980 3.940 ;
        RECT  0.160 3.285 0.420 3.940 ;
        RECT  0.000 3.440 0.160 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.785 0.925 4.885 1.185 ;
        RECT  4.785 2.175 4.885 2.775 ;
        RECT  4.625 0.925 4.785 3.100 ;
        RECT  1.340 2.940 4.625 3.100 ;
        RECT  3.705 0.925 3.865 2.755 ;
        RECT  3.605 0.925 3.705 1.185 ;
        RECT  3.605 2.155 3.705 2.755 ;
        RECT  1.785 2.595 3.605 2.755 ;
        RECT  2.910 1.430 3.010 1.690 ;
        RECT  2.750 0.945 2.910 2.400 ;
        RECT  2.585 0.945 2.750 1.205 ;
        RECT  2.555 2.240 2.750 2.400 ;
        RECT  1.785 0.935 1.820 1.195 ;
        RECT  1.625 0.935 1.785 2.755 ;
        RECT  1.560 0.935 1.625 1.195 ;
        RECT  1.520 2.115 1.625 2.755 ;
        RECT  1.340 1.410 1.445 1.685 ;
        RECT  1.330 1.410 1.340 3.100 ;
        RECT  1.180 0.925 1.330 3.100 ;
        RECT  1.170 0.925 1.180 2.630 ;
        RECT  0.820 0.925 1.170 1.085 ;
        RECT  0.820 2.395 1.170 2.630 ;
        RECT  0.560 0.825 0.820 1.085 ;
        RECT  0.560 2.180 0.820 2.780 ;
    END
END XOR2X2

MACRO XOR2X1
    CLASS CORE ;
    FOREIGN XOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 0.940 2.245 2.915 ;
        RECT  2.085 0.940 2.175 3.220 ;
        RECT  1.845 0.940 2.085 1.200 ;
        RECT  1.965 2.755 2.085 3.220 ;
        RECT  1.715 2.755 1.965 2.915 ;
        END
        ANTENNADIFFAREA     0.5382 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.125 1.290 1.255 1.580 ;
        RECT  0.965 1.290 1.125 1.890 ;
        RECT  0.830 1.630 0.965 1.890 ;
        END
        ANTENNAGATEAREA     0.1690 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 2.780 0.485 3.220 ;
        END
        ANTENNAGATEAREA     0.2340 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.090 -0.250 3.220 0.250 ;
        RECT  2.830 -0.250 3.090 0.405 ;
        RECT  1.060 -0.250 2.830 0.250 ;
        RECT  0.800 -0.250 1.060 1.110 ;
        RECT  0.000 -0.250 0.800 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.220 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.925 3.440 2.835 3.940 ;
        RECT  0.665 2.410 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.965 1.635 3.065 1.895 ;
        RECT  2.805 0.600 2.965 1.895 ;
        RECT  1.645 0.600 2.805 0.760 ;
        RECT  2.430 0.940 2.590 2.850 ;
        RECT  1.745 1.400 1.905 2.575 ;
        RECT  1.645 1.400 1.745 1.560 ;
        RECT  1.465 2.415 1.745 2.575 ;
        RECT  1.485 0.600 1.645 1.560 ;
        RECT  1.400 1.855 1.560 2.230 ;
        RECT  1.310 0.850 1.485 1.110 ;
        RECT  1.205 2.415 1.465 2.675 ;
        RECT  0.385 2.070 1.400 2.230 ;
        RECT  0.370 0.940 0.470 1.200 ;
        RECT  0.370 2.070 0.385 2.505 ;
        RECT  0.210 0.940 0.370 2.505 ;
        RECT  0.125 2.245 0.210 2.505 ;
    END
END XOR2X1

MACRO XOR2XL
    CLASS CORE ;
    FOREIGN XOR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.030 2.270 2.745 ;
        RECT  2.110 1.030 2.175 3.220 ;
        RECT  2.095 1.030 2.110 1.190 ;
        RECT  2.015 2.585 2.110 3.220 ;
        RECT  1.835 0.930 2.095 1.190 ;
        RECT  1.835 2.585 2.015 2.745 ;
        RECT  1.965 2.930 2.015 3.220 ;
        END
        ANTENNADIFFAREA     0.2377 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.465 1.090 1.725 ;
        RECT  0.585 1.290 0.795 1.725 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.790 0.500 3.140 ;
        RECT  0.125 2.790 0.335 3.220 ;
        RECT  0.120 2.790 0.125 3.140 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.220 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.955 -0.250 2.835 0.250 ;
        RECT  0.695 -0.250 0.955 1.110 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.220 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.955 3.440 2.835 3.940 ;
        RECT  0.695 2.335 0.955 3.940 ;
        RECT  0.000 3.440 0.695 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.805 0.590 2.965 1.735 ;
        RECT  1.580 0.590 2.805 0.750 ;
        RECT  2.455 0.930 2.615 2.705 ;
        RECT  1.770 1.400 1.930 2.405 ;
        RECT  1.580 1.400 1.770 1.560 ;
        RECT  1.525 2.245 1.770 2.405 ;
        RECT  1.430 1.785 1.590 2.065 ;
        RECT  1.420 0.590 1.580 1.560 ;
        RECT  1.265 2.245 1.525 2.595 ;
        RECT  0.385 1.905 1.430 2.065 ;
        RECT  1.265 0.930 1.420 1.190 ;
        RECT  0.285 0.915 0.385 1.175 ;
        RECT  0.285 1.905 0.385 2.485 ;
        RECT  0.125 0.915 0.285 2.485 ;
    END
END XOR2XL

MACRO CLKXOR2X8
    CLASS CORE ;
    FOREIGN CLKXOR2X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.015 1.000 9.075 2.760 ;
        RECT  8.755 1.000 9.015 3.020 ;
        RECT  8.675 1.000 8.755 2.760 ;
        RECT  8.405 1.000 8.675 2.420 ;
        RECT  7.445 1.000 8.405 1.400 ;
        RECT  7.995 2.020 8.405 2.420 ;
        RECT  7.735 2.020 7.995 3.190 ;
        END
        ANTENNADIFFAREA     1.3148 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.580 1.235 1.840 ;
        RECT  0.585 1.580 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.7020 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.795 1.565 2.055 1.825 ;
        RECT  1.715 1.665 1.795 1.825 ;
        RECT  1.505 1.665 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.7449 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.515 -0.250 9.660 0.250 ;
        RECT  9.255 -0.250 9.515 1.145 ;
        RECT  8.245 -0.250 9.255 0.250 ;
        RECT  7.985 -0.250 8.245 0.795 ;
        RECT  7.165 -0.250 7.985 0.250 ;
        RECT  6.905 -0.250 7.165 0.405 ;
        RECT  6.085 -0.250 6.905 0.250 ;
        RECT  5.825 -0.250 6.085 0.405 ;
        RECT  1.945 -0.250 5.825 0.250 ;
        RECT  1.685 -0.250 1.945 0.405 ;
        RECT  0.895 -0.250 1.685 0.250 ;
        RECT  0.635 -0.250 0.895 1.060 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.525 3.440 9.660 3.940 ;
        RECT  9.475 2.940 9.525 3.940 ;
        RECT  9.315 2.260 9.475 3.940 ;
        RECT  9.265 2.940 9.315 3.940 ;
        RECT  8.505 3.440 9.265 3.940 ;
        RECT  8.455 2.940 8.505 3.940 ;
        RECT  8.295 2.600 8.455 3.940 ;
        RECT  8.245 2.940 8.295 3.940 ;
        RECT  7.485 3.440 8.245 3.940 ;
        RECT  7.225 2.800 7.485 3.940 ;
        RECT  6.430 3.440 7.225 3.940 ;
        RECT  6.170 3.285 6.430 3.940 ;
        RECT  1.915 3.440 6.170 3.940 ;
        RECT  1.655 2.705 1.915 3.940 ;
        RECT  0.895 3.440 1.655 3.940 ;
        RECT  0.635 2.615 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.265 1.580 8.135 1.840 ;
        RECT  7.105 0.695 7.265 2.620 ;
        RECT  5.035 0.695 7.105 0.855 ;
        RECT  6.225 2.460 7.105 2.620 ;
        RECT  6.765 1.240 6.925 2.280 ;
        RECT  6.625 1.240 6.765 1.400 ;
        RECT  5.885 2.120 6.765 2.280 ;
        RECT  6.365 1.035 6.625 1.400 ;
        RECT  5.895 1.580 6.495 1.840 ;
        RECT  5.545 1.240 6.365 1.400 ;
        RECT  6.065 2.460 6.225 3.105 ;
        RECT  5.375 2.945 6.065 3.105 ;
        RECT  5.515 1.680 5.895 1.840 ;
        RECT  5.725 2.120 5.885 2.735 ;
        RECT  5.625 2.360 5.725 2.735 ;
        RECT  4.865 2.360 5.625 2.520 ;
        RECT  5.285 1.035 5.545 1.400 ;
        RECT  5.355 1.680 5.515 2.180 ;
        RECT  5.115 2.735 5.375 3.105 ;
        RECT  3.845 2.020 5.355 2.180 ;
        RECT  3.475 1.240 5.285 1.400 ;
        RECT  4.235 1.580 5.175 1.840 ;
        RECT  4.355 2.945 5.115 3.105 ;
        RECT  4.775 0.695 5.035 1.060 ;
        RECT  4.605 2.360 4.865 2.620 ;
        RECT  4.015 0.900 4.775 1.060 ;
        RECT  4.265 0.470 4.525 0.720 ;
        RECT  4.095 2.395 4.355 3.105 ;
        RECT  2.595 0.470 4.265 0.630 ;
        RECT  2.430 1.680 4.235 1.840 ;
        RECT  3.335 2.945 4.095 3.105 ;
        RECT  3.755 0.810 4.015 1.060 ;
        RECT  3.585 2.020 3.845 2.765 ;
        RECT  2.935 0.810 3.755 0.970 ;
        RECT  2.825 2.020 3.585 2.180 ;
        RECT  3.215 1.150 3.475 1.400 ;
        RECT  3.075 2.460 3.335 3.105 ;
        RECT  2.775 0.810 2.935 1.295 ;
        RECT  2.665 2.020 2.825 2.725 ;
        RECT  2.675 1.035 2.775 1.295 ;
        RECT  2.565 2.350 2.665 2.725 ;
        RECT  2.435 0.470 2.595 0.820 ;
        RECT  1.405 2.350 2.565 2.510 ;
        RECT  1.405 0.660 2.435 0.820 ;
        RECT  2.270 1.000 2.430 2.165 ;
        RECT  2.165 1.000 2.270 1.260 ;
        RECT  2.265 1.680 2.270 2.165 ;
        RECT  2.165 2.005 2.265 2.165 ;
        RECT  1.305 0.660 1.405 1.260 ;
        RECT  1.145 2.170 1.405 3.110 ;
        RECT  1.245 0.660 1.305 1.400 ;
        RECT  1.145 1.000 1.245 1.400 ;
        RECT  0.385 1.240 1.145 1.400 ;
        RECT  0.385 2.170 1.145 2.330 ;
        RECT  0.285 1.000 0.385 1.400 ;
        RECT  0.285 2.170 0.385 3.110 ;
        RECT  0.125 1.000 0.285 3.110 ;
    END
END CLKXOR2X8

MACRO CLKXOR2X4
    CLASS CORE ;
    FOREIGN CLKXOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.620 1.130 5.855 2.195 ;
        RECT  5.370 1.130 5.620 1.330 ;
        RECT  5.395 1.955 5.620 2.195 ;
        RECT  5.315 1.955 5.395 2.585 ;
        RECT  5.315 1.105 5.370 1.330 ;
        RECT  5.055 0.725 5.315 1.330 ;
        RECT  5.055 1.955 5.315 2.895 ;
        RECT  4.235 1.130 5.055 1.330 ;
        RECT  4.035 0.725 4.235 1.330 ;
        RECT  3.975 0.725 4.035 0.985 ;
        END
        ANTENNADIFFAREA     0.7924 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.585 0.385 1.845 ;
        RECT  0.125 1.585 0.335 2.400 ;
        END
        ANTENNAGATEAREA     0.3705 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.415 1.290 2.945 1.580 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.775 -0.250 5.980 0.250 ;
        RECT  4.515 -0.250 4.775 0.795 ;
        RECT  3.725 -0.250 4.515 0.250 ;
        RECT  3.465 -0.250 3.725 0.795 ;
        RECT  0.925 -0.250 3.465 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 3.440 5.980 3.940 ;
        RECT  5.595 2.555 5.855 3.940 ;
        RECT  4.805 3.440 5.595 3.940 ;
        RECT  4.545 2.595 4.805 3.940 ;
        RECT  1.325 3.440 4.545 3.940 ;
        RECT  1.065 3.285 1.325 3.940 ;
        RECT  0.385 3.440 1.065 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.030 1.510 5.290 1.770 ;
        RECT  4.875 1.610 5.030 1.770 ;
        RECT  4.715 1.610 4.875 2.305 ;
        RECT  3.255 2.145 4.715 2.305 ;
        RECT  4.035 1.645 4.295 1.965 ;
        RECT  3.285 1.805 4.035 1.965 ;
        RECT  3.770 3.000 4.030 3.260 ;
        RECT  3.765 3.000 3.770 3.160 ;
        RECT  3.505 2.630 3.765 3.160 ;
        RECT  0.945 2.925 3.505 3.085 ;
        RECT  3.125 0.820 3.285 1.965 ;
        RECT  2.995 2.145 3.255 2.745 ;
        RECT  3.065 0.820 3.125 0.980 ;
        RECT  2.745 1.805 3.125 1.965 ;
        RECT  2.805 0.720 3.065 0.980 ;
        RECT  2.235 2.440 2.995 2.600 ;
        RECT  2.585 1.805 2.745 2.260 ;
        RECT  2.485 2.000 2.585 2.260 ;
        RECT  2.295 0.720 2.555 1.110 ;
        RECT  2.235 0.950 2.295 1.110 ;
        RECT  2.075 0.950 2.235 2.600 ;
        RECT  1.975 2.000 2.075 2.600 ;
        RECT  1.785 0.510 2.045 0.770 ;
        RECT  1.495 1.265 1.895 1.525 ;
        RECT  0.385 0.610 1.785 0.770 ;
        RECT  1.465 1.955 1.725 2.215 ;
        RECT  1.395 1.035 1.495 1.525 ;
        RECT  1.395 1.955 1.465 2.115 ;
        RECT  1.235 1.035 1.395 2.115 ;
        RECT  0.785 1.245 0.945 3.085 ;
        RECT  0.385 1.245 0.785 1.405 ;
        RECT  0.525 2.135 0.785 2.735 ;
        RECT  0.125 0.610 0.385 1.405 ;
    END
END CLKXOR2X4

MACRO CLKXOR2X2
    CLASS CORE ;
    FOREIGN CLKXOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.545 0.880 3.555 1.170 ;
        RECT  3.545 2.745 3.555 2.995 ;
        RECT  3.490 0.880 3.545 2.995 ;
        RECT  3.385 0.880 3.490 3.195 ;
        RECT  3.370 0.880 3.385 1.355 ;
        RECT  3.230 2.595 3.385 3.195 ;
        RECT  3.345 0.880 3.370 1.295 ;
        RECT  3.285 1.035 3.345 1.295 ;
        END
        ANTENNADIFFAREA     0.6017 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.860 1.020 1.020 2.270 ;
        RECT  0.795 2.110 0.860 2.270 ;
        RECT  0.585 2.110 0.795 2.400 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.095 0.340 1.590 ;
        END
        ANTENNAGATEAREA     0.2184 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 -0.250 3.680 0.250 ;
        RECT  2.690 -0.250 2.950 0.405 ;
        RECT  0.815 -0.250 2.690 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 3.440 3.680 3.940 ;
        RECT  2.690 2.945 2.950 3.940 ;
        RECT  0.850 3.440 2.690 3.940 ;
        RECT  0.590 3.285 0.850 3.940 ;
        RECT  0.000 3.440 0.590 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.020 1.585 3.180 2.400 ;
        RECT  2.840 2.240 3.020 2.400 ;
        RECT  2.680 0.585 2.840 1.960 ;
        RECT  2.680 2.240 2.840 2.740 ;
        RECT  2.085 0.585 2.680 0.745 ;
        RECT  2.670 1.800 2.680 1.960 ;
        RECT  1.960 2.580 2.680 2.740 ;
        RECT  2.510 1.800 2.670 2.060 ;
        RECT  2.340 1.035 2.500 1.610 ;
        RECT  2.310 2.240 2.410 2.400 ;
        RECT  2.310 1.450 2.340 1.610 ;
        RECT  2.150 1.450 2.310 2.400 ;
        RECT  1.435 3.100 2.240 3.260 ;
        RECT  1.925 0.585 2.085 0.930 ;
        RECT  1.900 1.110 1.960 2.740 ;
        RECT  1.510 0.770 1.925 0.930 ;
        RECT  1.800 1.110 1.900 2.780 ;
        RECT  1.640 2.180 1.800 2.780 ;
        RECT  1.155 0.430 1.640 0.590 ;
        RECT  1.390 0.770 1.510 1.135 ;
        RECT  1.275 2.945 1.435 3.260 ;
        RECT  1.350 0.770 1.390 2.710 ;
        RECT  1.230 0.925 1.350 2.710 ;
        RECT  0.385 2.945 1.275 3.105 ;
        RECT  1.130 2.450 1.230 2.710 ;
        RECT  0.995 0.430 1.155 0.745 ;
        RECT  0.680 0.585 0.995 0.745 ;
        RECT  0.520 0.585 0.680 1.930 ;
        RECT  0.125 0.755 0.520 0.915 ;
        RECT  0.385 1.770 0.520 1.930 ;
        RECT  0.225 1.770 0.385 3.105 ;
        RECT  0.125 2.280 0.225 2.540 ;
    END
END CLKXOR2X2

MACRO CLKXOR2X1
    CLASS CORE ;
    FOREIGN CLKXOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.545 0.880 3.555 2.585 ;
        RECT  3.345 0.880 3.545 2.615 ;
        RECT  3.335 0.945 3.345 1.295 ;
        RECT  3.285 2.355 3.345 2.615 ;
        RECT  3.285 1.035 3.335 1.295 ;
        END
        ANTENNADIFFAREA     0.3196 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 1.115 1.105 2.270 ;
        RECT  0.905 1.910 0.945 2.270 ;
        RECT  0.795 2.110 0.905 2.270 ;
        RECT  0.585 2.110 0.795 2.400 ;
        END
        ANTENNAGATEAREA     0.0949 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.170 0.385 1.590 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.965 -0.250 3.680 0.250 ;
        RECT  2.705 -0.250 2.965 0.405 ;
        RECT  0.955 -0.250 2.705 0.250 ;
        RECT  0.695 -0.250 0.955 0.650 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 3.440 3.680 3.940 ;
        RECT  2.710 2.945 2.970 3.940 ;
        RECT  0.850 3.440 2.710 3.940 ;
        RECT  0.590 3.285 0.850 3.940 ;
        RECT  0.000 3.440 0.590 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.060 1.820 3.160 2.080 ;
        RECT  2.900 1.820 3.060 2.740 ;
        RECT  2.795 0.585 2.955 1.635 ;
        RECT  1.795 2.580 2.900 2.740 ;
        RECT  1.535 0.585 2.795 0.745 ;
        RECT  2.720 1.475 2.795 1.635 ;
        RECT  2.560 1.475 2.720 1.985 ;
        RECT  2.315 1.725 2.560 1.985 ;
        RECT  2.380 1.035 2.535 1.295 ;
        RECT  2.135 2.240 2.390 2.400 ;
        RECT  2.220 1.035 2.380 1.540 ;
        RECT  2.135 1.380 2.220 1.540 ;
        RECT  1.975 1.380 2.135 2.400 ;
        RECT  1.725 2.920 1.985 3.180 ;
        RECT  1.795 0.960 1.965 1.120 ;
        RECT  1.635 0.960 1.795 2.740 ;
        RECT  0.385 2.920 1.725 3.080 ;
        RECT  1.455 0.450 1.535 0.745 ;
        RECT  1.295 0.450 1.455 2.710 ;
        RECT  1.275 0.450 1.295 0.610 ;
        RECT  1.075 2.450 1.295 2.710 ;
        RECT  0.565 0.830 0.725 1.930 ;
        RECT  0.385 0.830 0.565 0.990 ;
        RECT  0.385 1.770 0.565 1.930 ;
        RECT  0.125 0.730 0.385 0.990 ;
        RECT  0.225 1.770 0.385 3.080 ;
        RECT  0.125 2.280 0.225 2.540 ;
    END
END CLKXOR2X1

MACRO OA22X4
    CLASS CORE ;
    FOREIGN OA22X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.700 4.015 2.400 ;
        RECT  3.805 1.315 4.005 2.710 ;
        RECT  3.555 1.315 3.805 1.515 ;
        RECT  3.295 2.510 3.805 2.710 ;
        RECT  3.505 1.105 3.555 1.515 ;
        RECT  3.305 0.635 3.505 1.515 ;
        RECT  3.245 0.635 3.305 1.235 ;
        RECT  3.035 2.510 3.295 3.195 ;
        END
        ANTENNADIFFAREA     0.7486 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.290 2.770 1.960 ;
        END
        ANTENNAGATEAREA     0.2561 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.175 1.990 ;
        RECT  1.815 1.290 1.965 1.930 ;
        END
        ANTENNAGATEAREA     0.2561 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.525 1.695 0.625 1.955 ;
        RECT  0.365 1.695 0.525 2.270 ;
        RECT  0.335 2.110 0.365 2.270 ;
        RECT  0.125 2.110 0.335 2.400 ;
        END
        ANTENNAGATEAREA     0.2561 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 2.110 1.715 2.400 ;
        RECT  1.405 1.700 1.635 2.400 ;
        RECT  1.330 1.700 1.405 1.960 ;
        END
        ANTENNAGATEAREA     0.2561 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 -0.250 4.140 0.250 ;
        RECT  3.755 -0.250 4.015 1.120 ;
        RECT  2.995 -0.250 3.755 0.250 ;
        RECT  2.735 -0.250 2.995 1.070 ;
        RECT  1.975 -0.250 2.735 0.250 ;
        RECT  1.715 -0.250 1.975 0.760 ;
        RECT  0.000 -0.250 1.715 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.835 3.440 4.140 3.940 ;
        RECT  3.575 2.935 3.835 3.940 ;
        RECT  2.755 3.440 3.575 3.940 ;
        RECT  2.495 2.595 2.755 3.940 ;
        RECT  0.885 3.440 2.495 3.940 ;
        RECT  0.625 2.545 0.885 3.940 ;
        RECT  0.000 3.440 0.625 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.215 1.695 3.335 1.955 ;
        RECT  3.055 1.695 3.215 2.330 ;
        RECT  2.055 2.170 3.055 2.330 ;
        RECT  2.385 0.665 2.485 0.925 ;
        RECT  2.225 0.665 2.385 1.110 ;
        RECT  1.455 0.950 2.225 1.110 ;
        RECT  1.905 2.170 2.055 2.740 ;
        RECT  1.895 2.170 1.905 3.180 ;
        RECT  1.645 2.580 1.895 3.180 ;
        RECT  1.225 2.580 1.645 2.740 ;
        RECT  1.195 0.650 1.455 1.320 ;
        RECT  1.065 2.140 1.225 2.740 ;
        RECT  0.435 0.650 1.195 0.810 ;
        RECT  0.965 2.140 1.065 2.300 ;
        RECT  0.805 0.990 0.965 2.300 ;
        RECT  0.685 0.990 0.805 1.250 ;
        RECT  0.175 0.650 0.435 1.250 ;
    END
END OA22X4

MACRO OA22X2
    CLASS CORE ;
    FOREIGN OA22X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 0.695 3.095 2.995 ;
        RECT  2.935 0.695 2.975 3.195 ;
        RECT  2.835 0.695 2.935 1.295 ;
        RECT  2.885 2.110 2.935 3.195 ;
        RECT  2.715 2.595 2.885 3.195 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.475 2.175 1.990 ;
        RECT  1.895 1.475 1.965 1.985 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.475 1.715 1.990 ;
        RECT  1.285 1.475 1.505 1.735 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.310 0.335 2.365 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.110 1.255 2.400 ;
        RECT  0.945 1.475 1.105 2.400 ;
        RECT  0.855 1.475 0.945 1.735 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 -0.250 3.220 0.250 ;
        RECT  1.835 -0.250 2.545 0.405 ;
        RECT  0.000 -0.250 1.835 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.435 3.440 3.220 3.940 ;
        RECT  2.175 2.605 2.435 3.940 ;
        RECT  1.835 2.605 2.175 2.765 ;
        RECT  0.385 3.440 2.175 3.940 ;
        RECT  0.125 2.545 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.705 1.585 2.755 1.845 ;
        RECT  2.595 1.585 2.705 2.400 ;
        RECT  2.545 1.590 2.595 2.400 ;
        RECT  1.595 2.240 2.545 2.400 ;
        RECT  1.895 1.035 2.155 1.295 ;
        RECT  1.245 1.035 1.895 1.195 ;
        RECT  1.435 2.240 1.595 2.740 ;
        RECT  1.235 2.580 1.435 2.740 ;
        RECT  1.085 0.435 1.245 1.195 ;
        RECT  0.975 2.580 1.235 2.840 ;
        RECT  0.985 0.435 1.085 0.595 ;
        RECT  0.765 2.580 0.975 2.740 ;
        RECT  0.675 0.985 0.785 1.245 ;
        RECT  0.675 2.205 0.765 2.740 ;
        RECT  0.605 0.985 0.675 2.740 ;
        RECT  0.515 0.985 0.605 2.365 ;
    END
END OA22X2

MACRO OA22X1
    CLASS CORE ;
    FOREIGN OA22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.830 2.660 2.995 ;
        RECT  2.625 0.735 2.635 2.995 ;
        RECT  2.500 0.735 2.625 3.215 ;
        RECT  2.425 0.735 2.500 1.990 ;
        RECT  2.465 2.610 2.500 3.215 ;
        RECT  2.345 2.955 2.465 3.215 ;
        RECT  2.375 0.735 2.425 0.995 ;
        END
        ANTENNADIFFAREA     0.3366 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.110 1.945 2.400 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.670 1.410 1.930 ;
        RECT  0.980 1.670 1.330 1.990 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.105 0.400 1.590 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 2.175 1.070 2.435 ;
        RECT  0.585 2.110 0.795 2.435 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.070 -0.250 2.760 0.250 ;
        RECT  1.810 -0.250 2.070 1.150 ;
        RECT  0.000 -0.250 1.810 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.095 3.440 2.760 3.940 ;
        RECT  1.835 2.955 2.095 3.940 ;
        RECT  0.390 3.440 1.835 3.940 ;
        RECT  0.130 2.955 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.285 2.170 2.320 2.430 ;
        RECT  2.125 2.170 2.285 2.775 ;
        RECT  1.240 2.615 2.125 2.775 ;
        RECT  2.000 1.625 2.100 1.885 ;
        RECT  1.840 1.330 2.000 1.885 ;
        RECT  1.470 1.330 1.840 1.490 ;
        RECT  1.370 0.735 1.470 1.490 ;
        RECT  1.310 0.570 1.370 1.490 ;
        RECT  1.210 0.570 1.310 0.995 ;
        RECT  0.980 2.615 1.240 2.995 ;
        RECT  0.385 0.570 1.210 0.730 ;
        RECT  0.405 2.615 0.980 2.775 ;
        RECT  0.800 0.960 0.900 1.220 ;
        RECT  0.640 0.960 0.800 1.930 ;
        RECT  0.405 1.770 0.640 1.930 ;
        RECT  0.245 1.770 0.405 2.775 ;
        RECT  0.125 0.470 0.385 0.730 ;
    END
END OA22X1

MACRO OA22XL
    CLASS CORE ;
    FOREIGN OA22XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 2.245 2.670 3.215 ;
        RECT  2.510 0.735 2.635 3.215 ;
        RECT  2.475 0.735 2.510 2.405 ;
        RECT  2.345 2.955 2.510 3.215 ;
        RECT  2.425 0.735 2.475 2.175 ;
        RECT  2.375 0.735 2.425 0.995 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.890 2.110 2.175 2.400 ;
        RECT  1.630 2.065 1.890 2.400 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.670 1.410 1.990 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.105 0.400 1.590 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 2.175 1.070 2.435 ;
        RECT  0.585 2.110 0.795 2.435 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.050 -0.250 2.760 0.250 ;
        RECT  1.790 -0.250 2.050 1.150 ;
        RECT  0.000 -0.250 1.790 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.095 3.440 2.760 3.940 ;
        RECT  1.835 2.955 2.095 3.940 ;
        RECT  0.390 3.440 1.835 3.940 ;
        RECT  0.130 2.955 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.070 2.595 2.330 2.775 ;
        RECT  2.000 1.625 2.100 1.885 ;
        RECT  1.240 2.615 2.070 2.775 ;
        RECT  1.840 1.330 2.000 1.885 ;
        RECT  1.470 1.330 1.840 1.490 ;
        RECT  1.370 0.735 1.470 1.490 ;
        RECT  1.310 0.580 1.370 1.490 ;
        RECT  1.210 0.580 1.310 0.995 ;
        RECT  0.980 2.615 1.240 2.995 ;
        RECT  0.385 0.580 1.210 0.740 ;
        RECT  0.405 2.615 0.980 2.775 ;
        RECT  0.800 0.970 0.900 1.230 ;
        RECT  0.640 0.970 0.800 1.930 ;
        RECT  0.405 1.770 0.640 1.930 ;
        RECT  0.245 1.770 0.405 2.775 ;
        RECT  0.125 0.480 0.385 0.740 ;
    END
END OA22XL

MACRO OA21X4
    CLASS CORE ;
    FOREIGN OA21X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.675 0.535 2.935 3.045 ;
        RECT  2.425 1.700 2.675 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.690 1.700 1.715 1.990 ;
        RECT  1.505 1.635 1.690 1.990 ;
        RECT  1.285 1.635 1.505 1.930 ;
        END
        ANTENNAGATEAREA     0.2405 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.505 0.375 1.990 ;
        END
        ANTENNAGATEAREA     0.2795 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.690 1.580 1.015 1.990 ;
        RECT  0.585 1.700 0.690 1.990 ;
        END
        ANTENNAGATEAREA     0.2795 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.475 -0.250 3.680 0.250 ;
        RECT  3.215 -0.250 3.475 1.175 ;
        RECT  2.425 -0.250 3.215 0.250 ;
        RECT  2.165 -0.250 2.425 1.095 ;
        RECT  0.895 -0.250 2.165 0.250 ;
        RECT  0.635 -0.250 0.895 0.900 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.475 3.440 3.680 3.940 ;
        RECT  3.215 2.215 3.475 3.940 ;
        RECT  2.185 3.440 3.215 3.940 ;
        RECT  1.925 2.555 2.185 3.940 ;
        RECT  0.385 3.440 1.925 3.940 ;
        RECT  0.125 2.200 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.060 1.585 2.155 1.845 ;
        RECT  2.055 1.295 2.060 1.845 ;
        RECT  1.915 1.295 2.055 2.360 ;
        RECT  1.895 0.695 1.915 2.360 ;
        RECT  1.655 0.695 1.895 1.455 ;
        RECT  1.235 2.200 1.895 2.360 ;
        RECT  1.145 0.695 1.405 1.295 ;
        RECT  0.975 2.200 1.235 2.800 ;
        RECT  0.385 1.135 1.145 1.295 ;
        RECT  0.125 0.695 0.385 1.295 ;
    END
END OA21X4

MACRO OA21X2
    CLASS CORE ;
    FOREIGN OA21X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 0.745 2.635 2.170 ;
        RECT  2.180 0.745 2.425 1.005 ;
        RECT  2.175 2.010 2.425 2.170 ;
        RECT  2.120 2.010 2.175 2.995 ;
        RECT  1.960 2.010 2.120 3.125 ;
        RECT  1.835 2.525 1.960 3.125 ;
        END
        ANTENNADIFFAREA     0.4726 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.340 1.725 1.440 1.985 ;
        RECT  1.180 0.880 1.340 1.985 ;
        RECT  1.045 0.880 1.180 1.170 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.375 1.990 ;
        RECT  0.115 1.510 0.125 1.770 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.615 0.910 2.005 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 -0.250 2.760 0.250 ;
        RECT  1.760 -0.250 2.360 0.405 ;
        RECT  0.845 -0.250 1.760 0.250 ;
        RECT  0.585 -0.250 0.845 1.270 ;
        RECT  0.000 -0.250 0.585 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 3.440 2.760 3.940 ;
        RECT  2.375 2.525 2.635 3.940 ;
        RECT  1.550 3.440 2.375 3.940 ;
        RECT  1.290 3.285 1.550 3.940 ;
        RECT  0.385 3.440 1.290 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.985 1.210 2.245 1.830 ;
        RECT  1.610 1.210 1.985 1.470 ;
        RECT  1.780 1.670 1.985 1.830 ;
        RECT  1.620 1.670 1.780 2.345 ;
        RECT  1.130 2.185 1.620 2.345 ;
        RECT  0.970 2.185 1.130 2.725 ;
        RECT  0.870 2.465 0.970 2.725 ;
    END
END OA21X2

MACRO OA21X1
    CLASS CORE ;
    FOREIGN OA21X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.450 2.110 2.635 2.400 ;
        RECT  2.430 2.110 2.450 2.555 ;
        RECT  2.270 1.030 2.430 2.555 ;
        RECT  2.110 1.030 2.270 1.290 ;
        RECT  2.110 1.955 2.270 2.555 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 1.405 1.545 1.665 ;
        RECT  1.285 1.010 1.445 1.665 ;
        RECT  1.255 1.010 1.285 1.170 ;
        RECT  1.045 0.880 1.255 1.170 ;
        END
        ANTENNAGATEAREA     0.0611 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.115 1.510 0.375 1.990 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.600 1.015 1.990 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 -0.250 2.760 0.250 ;
        RECT  2.110 -0.250 2.370 0.780 ;
        RECT  0.835 -0.250 2.110 0.250 ;
        RECT  0.575 -0.250 0.835 1.295 ;
        RECT  0.000 -0.250 0.575 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 3.440 2.760 3.940 ;
        RECT  1.565 2.190 1.825 3.940 ;
        RECT  0.415 3.440 1.565 3.940 ;
        RECT  0.155 2.170 0.415 3.940 ;
        RECT  0.000 3.440 0.155 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.895 1.485 2.075 1.745 ;
        RECT  1.735 0.490 1.895 2.010 ;
        RECT  1.550 0.490 1.735 0.750 ;
        RECT  1.385 1.850 1.735 2.010 ;
        RECT  1.235 1.850 1.385 2.390 ;
        RECT  1.225 1.850 1.235 2.430 ;
        RECT  0.975 2.170 1.225 2.430 ;
    END
END OA21X1

MACRO OA21XL
    CLASS CORE ;
    FOREIGN OA21XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.310 2.210 2.250 ;
        RECT  2.050 0.440 2.175 2.400 ;
        RECT  1.915 0.440 2.050 1.470 ;
        RECT  1.965 2.090 2.050 2.400 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 1.575 1.380 1.835 ;
        RECT  1.105 0.880 1.265 1.835 ;
        RECT  1.045 0.880 1.105 1.170 ;
        END
        ANTENNAGATEAREA     0.0572 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.510 0.400 1.990 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.505 0.925 1.990 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.605 -0.250 2.300 0.250 ;
        RECT  1.345 -0.250 1.605 0.405 ;
        RECT  0.580 -0.250 1.345 0.250 ;
        RECT  0.320 -0.250 0.580 1.125 ;
        RECT  0.000 -0.250 0.320 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 3.440 2.300 3.940 ;
        RECT  1.375 2.680 1.635 3.940 ;
        RECT  0.385 3.440 1.375 3.940 ;
        RECT  0.125 2.750 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.720 1.650 1.870 1.910 ;
        RECT  1.560 1.045 1.720 2.330 ;
        RECT  1.445 1.045 1.560 1.305 ;
        RECT  1.095 2.170 1.560 2.330 ;
        RECT  0.835 2.170 1.095 2.430 ;
    END
END OA21XL

MACRO OAI2BB2X4
    CLASS CORE ;
    FOREIGN OAI2BB2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.305 1.515 6.315 3.080 ;
        RECT  6.105 0.975 6.305 3.080 ;
        RECT  5.110 0.975 6.105 1.175 ;
        RECT  6.055 2.140 6.105 3.080 ;
        RECT  4.895 2.710 6.055 2.910 ;
        RECT  4.910 0.975 5.110 1.475 ;
        RECT  4.190 1.275 4.910 1.475 ;
        RECT  4.635 2.710 4.895 2.970 ;
        RECT  3.815 2.710 4.635 2.910 ;
        RECT  3.990 0.810 4.190 1.475 ;
        RECT  3.920 0.810 3.990 1.410 ;
        RECT  3.555 2.710 3.815 2.970 ;
        RECT  2.410 2.710 3.555 2.910 ;
        RECT  2.150 2.585 2.410 3.185 ;
        END
        ANTENNADIFFAREA     1.7285 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.930 1.710 5.030 1.970 ;
        RECT  4.770 1.710 4.930 2.190 ;
        RECT  4.725 1.925 4.770 2.190 ;
        RECT  3.190 2.030 4.725 2.190 ;
        RECT  3.090 1.745 3.190 2.190 ;
        RECT  2.930 1.455 3.090 2.190 ;
        RECT  1.750 1.455 2.930 1.615 ;
        RECT  1.540 1.455 1.750 1.990 ;
        RECT  1.490 1.460 1.540 1.990 ;
        END
        ANTENNAGATEAREA     0.7358 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.660 1.385 5.920 1.645 ;
        RECT  5.500 1.485 5.660 1.645 ;
        RECT  5.340 1.485 5.500 2.530 ;
        RECT  5.210 2.335 5.340 2.530 ;
        RECT  2.750 2.370 5.210 2.530 ;
        RECT  2.590 1.795 2.750 2.530 ;
        RECT  2.425 1.795 2.590 2.175 ;
        RECT  2.175 1.795 2.425 1.995 ;
        RECT  1.970 1.795 2.175 2.400 ;
        RECT  1.965 1.800 1.970 2.400 ;
        END
        ANTENNAGATEAREA     0.7358 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.555 1.280 2.025 ;
        END
        ANTENNAGATEAREA     0.2587 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.445 0.485 1.990 ;
        END
        ANTENNAGATEAREA     0.2587 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 -0.250 6.440 0.250 ;
        RECT  6.055 -0.250 6.315 0.795 ;
        RECT  5.230 -0.250 6.055 0.250 ;
        RECT  4.970 -0.250 5.230 0.405 ;
        RECT  3.130 -0.250 4.970 0.250 ;
        RECT  2.870 -0.250 3.130 0.405 ;
        RECT  1.605 -0.250 2.870 0.250 ;
        RECT  1.345 -0.250 1.605 0.735 ;
        RECT  0.385 -0.250 1.345 0.250 ;
        RECT  0.125 -0.250 0.385 1.080 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.460 3.440 6.440 3.940 ;
        RECT  5.200 3.285 5.460 3.940 ;
        RECT  4.355 3.440 5.200 3.940 ;
        RECT  4.095 3.285 4.355 3.940 ;
        RECT  3.275 3.440 4.095 3.940 ;
        RECT  3.015 3.285 3.275 3.940 ;
        RECT  1.505 3.440 3.015 3.940 ;
        RECT  1.245 2.210 1.505 3.940 ;
        RECT  0.385 3.440 1.245 3.940 ;
        RECT  0.125 2.215 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.510 0.500 5.770 0.760 ;
        RECT  4.690 0.600 5.510 0.760 ;
        RECT  4.430 0.470 4.690 1.095 ;
        RECT  3.670 0.470 4.430 0.630 ;
        RECT  3.615 1.590 3.810 1.850 ;
        RECT  3.410 0.470 3.670 0.935 ;
        RECT  3.455 1.115 3.615 1.850 ;
        RECT  1.205 1.115 3.455 1.275 ;
        RECT  2.115 0.775 3.410 0.935 ;
        RECT  1.855 0.680 2.115 0.935 ;
        RECT  0.945 1.035 1.205 1.295 ;
        RECT  0.825 1.135 0.945 1.295 ;
        RECT  0.825 2.220 0.925 2.820 ;
        RECT  0.665 1.135 0.825 2.820 ;
    END
END OAI2BB2X4

MACRO OAI2BB2X2
    CLASS CORE ;
    FOREIGN OAI2BB2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.335 1.215 4.495 2.445 ;
        RECT  4.015 1.215 4.335 1.375 ;
        RECT  4.265 2.110 4.335 2.445 ;
        RECT  3.715 2.285 4.265 2.445 ;
        RECT  3.855 0.925 4.015 1.375 ;
        RECT  2.985 0.925 3.855 1.085 ;
        RECT  3.455 2.285 3.715 2.885 ;
        RECT  2.635 2.285 3.455 2.445 ;
        RECT  2.725 0.820 2.985 1.085 ;
        RECT  2.515 2.285 2.635 2.585 ;
        RECT  2.450 2.285 2.515 2.740 ;
        RECT  2.355 2.285 2.450 2.840 ;
        RECT  2.055 2.580 2.355 2.840 ;
        END
        ANTENNADIFFAREA     0.9748 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 1.265 3.640 1.425 ;
        RECT  3.380 1.265 3.540 1.765 ;
        RECT  3.345 1.515 3.380 1.765 ;
        RECT  1.715 1.605 3.345 1.765 ;
        RECT  1.440 1.605 1.715 2.105 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.055 1.555 4.155 1.815 ;
        RECT  3.895 1.555 4.055 2.105 ;
        RECT  3.830 1.925 3.895 2.105 ;
        RECT  2.175 1.945 3.830 2.105 ;
        RECT  1.965 1.945 2.175 2.400 ;
        RECT  1.920 1.945 1.965 2.105 ;
        END
        ANTENNAGATEAREA     0.3640 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.010 1.545 1.255 2.070 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.120 1.465 0.395 1.990 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 -0.250 4.600 0.250 ;
        RECT  3.815 -0.250 4.075 0.405 ;
        RECT  2.075 -0.250 3.815 0.250 ;
        RECT  1.815 -0.250 2.075 0.405 ;
        RECT  0.385 -0.250 1.815 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.175 3.440 4.600 3.940 ;
        RECT  2.915 2.725 3.175 3.940 ;
        RECT  1.465 3.440 2.915 3.940 ;
        RECT  1.205 2.515 1.465 3.940 ;
        RECT  0.385 3.440 1.205 3.940 ;
        RECT  0.125 2.215 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.375 0.775 4.475 1.035 ;
        RECT  4.215 0.585 4.375 1.035 ;
        RECT  3.495 0.585 4.215 0.745 ;
        RECT  3.230 0.480 3.495 0.745 ;
        RECT  2.475 0.480 3.230 0.640 ;
        RECT  1.850 1.265 3.140 1.425 ;
        RECT  2.315 0.480 2.475 1.035 ;
        RECT  2.215 0.625 2.315 1.035 ;
        RECT  1.495 0.625 2.215 0.785 ;
        RECT  1.690 1.165 1.850 1.425 ;
        RECT  1.095 1.165 1.690 1.325 ;
        RECT  1.235 0.525 1.495 0.785 ;
        RECT  0.835 1.035 1.095 1.325 ;
        RECT  0.825 2.260 0.925 2.520 ;
        RECT  0.825 1.165 0.835 1.325 ;
        RECT  0.665 1.165 0.825 2.520 ;
    END
END OAI2BB2X2

MACRO OAI2BB2X1
    CLASS CORE ;
    FOREIGN OAI2BB2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.985 1.105 3.095 2.400 ;
        RECT  2.825 0.845 2.985 2.670 ;
        RECT  2.725 0.845 2.825 1.105 ;
        RECT  2.060 2.510 2.825 2.670 ;
        END
        ANTENNADIFFAREA     0.4911 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.450 1.230 1.715 1.730 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.355 2.180 1.990 ;
        RECT  1.965 1.290 2.175 1.990 ;
        RECT  1.920 1.730 1.965 1.990 ;
        END
        ANTENNAGATEAREA     0.1820 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.010 1.480 1.255 1.990 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.235 1.570 0.485 2.000 ;
        RECT  0.125 1.700 0.235 2.000 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.075 -0.250 3.220 0.250 ;
        RECT  1.815 -0.250 2.075 0.405 ;
        RECT  0.385 -0.250 1.815 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.865 3.440 3.220 3.940 ;
        RECT  2.605 2.920 2.865 3.940 ;
        RECT  1.465 3.440 2.605 3.940 ;
        RECT  1.205 2.515 1.465 3.940 ;
        RECT  0.385 3.440 1.205 3.940 ;
        RECT  0.125 2.215 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.485 1.715 2.645 2.330 ;
        RECT  0.830 2.170 2.485 2.330 ;
        RECT  2.375 0.835 2.475 1.095 ;
        RECT  2.215 0.625 2.375 1.095 ;
        RECT  1.485 0.625 2.215 0.785 ;
        RECT  1.225 0.525 1.485 0.785 ;
        RECT  0.865 1.035 1.125 1.295 ;
        RECT  0.830 1.085 0.865 1.295 ;
        RECT  0.665 1.085 0.830 2.330 ;
    END
END OAI2BB2X1

MACRO OAI2BB2XL
    CLASS CORE ;
    FOREIGN OAI2BB2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 0.790 2.640 2.745 ;
        RECT  2.480 0.790 2.635 2.810 ;
        RECT  2.425 0.790 2.480 1.355 ;
        RECT  2.425 2.515 2.480 2.810 ;
        RECT  2.360 0.790 2.425 1.050 ;
        RECT  1.900 2.515 2.425 2.675 ;
        END
        ANTENNADIFFAREA     0.2599 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.700 1.715 1.990 ;
        RECT  1.240 1.710 1.505 1.970 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.175 1.580 ;
        RECT  1.820 1.290 1.965 1.490 ;
        RECT  1.560 1.230 1.820 1.490 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 2.520 1.040 2.810 ;
        END
        ANTENNAGATEAREA     0.0572 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.465 0.445 1.990 ;
        END
        ANTENNAGATEAREA     0.0572 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.710 -0.250 2.760 0.250 ;
        RECT  1.450 -0.250 1.710 0.405 ;
        RECT  0.385 -0.250 1.450 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 3.440 2.760 3.940 ;
        RECT  2.300 3.285 2.560 3.940 ;
        RECT  1.440 3.440 2.300 3.940 ;
        RECT  1.180 3.285 1.440 3.940 ;
        RECT  0.385 3.440 1.180 3.940 ;
        RECT  0.125 2.860 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.040 1.925 2.300 2.335 ;
        RECT  2.010 0.780 2.110 1.040 ;
        RECT  1.030 2.175 2.040 2.335 ;
        RECT  1.850 0.625 2.010 1.040 ;
        RECT  1.140 0.625 1.850 0.785 ;
        RECT  0.880 0.525 1.140 0.785 ;
        RECT  1.030 1.035 1.125 1.295 ;
        RECT  0.865 1.035 1.030 2.335 ;
        RECT  0.555 2.175 0.865 2.335 ;
    END
END OAI2BB2XL

MACRO OAI2BB1X4
    CLASS CORE ;
    FOREIGN OAI2BB1X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 0.470 4.015 2.585 ;
        RECT  3.740 0.470 3.805 1.170 ;
        RECT  3.475 2.345 3.805 2.585 ;
        RECT  2.450 0.915 3.740 1.115 ;
        RECT  3.215 2.345 3.475 2.970 ;
        RECT  2.455 2.345 3.215 2.545 ;
        RECT  2.195 2.345 2.455 2.970 ;
        RECT  2.100 0.800 2.450 1.115 ;
        END
        ANTENNADIFFAREA     1.4700 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.810 1.295 3.070 1.710 ;
        RECT  1.715 1.295 2.810 1.455 ;
        RECT  1.655 0.880 1.715 1.455 ;
        RECT  1.495 0.880 1.655 1.665 ;
        END
        ANTENNAGATEAREA     0.5928 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.470 0.345 2.055 ;
        END
        ANTENNAGATEAREA     0.2548 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.290 1.255 1.580 ;
        RECT  0.865 1.290 1.230 1.825 ;
        END
        ANTENNAGATEAREA     0.2548 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.180 -0.250 4.140 0.250 ;
        RECT  2.920 -0.250 3.180 0.705 ;
        RECT  1.205 -0.250 2.920 0.250 ;
        RECT  0.945 -0.250 1.205 1.075 ;
        RECT  0.000 -0.250 0.945 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.845 4.015 3.940 ;
        RECT  2.965 3.440 3.755 3.940 ;
        RECT  2.705 2.785 2.965 3.940 ;
        RECT  1.740 3.440 2.705 3.940 ;
        RECT  1.480 2.395 1.740 3.940 ;
        RECT  0.450 3.440 1.480 3.940 ;
        RECT  0.190 2.530 0.450 3.940 ;
        RECT  0.000 3.440 0.190 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.405 1.575 3.565 2.165 ;
        RECT  2.190 2.005 3.405 2.165 ;
        RECT  1.930 1.635 2.190 2.165 ;
        RECT  1.045 2.005 1.930 2.165 ;
        RECT  0.785 2.005 1.045 3.015 ;
        RECT  0.685 2.005 0.785 2.165 ;
        RECT  0.525 1.125 0.685 2.165 ;
        RECT  0.385 1.125 0.525 1.285 ;
        RECT  0.125 0.585 0.385 1.285 ;
    END
END OAI2BB1X4

MACRO OAI2BB1X2
    CLASS CORE ;
    FOREIGN OAI2BB1X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 0.930 3.095 2.275 ;
        RECT  2.115 0.930 2.935 1.090 ;
        RECT  2.175 2.115 2.935 2.275 ;
        RECT  2.130 2.110 2.175 2.995 ;
        RECT  1.965 2.110 2.130 3.205 ;
        RECT  1.855 0.830 2.115 1.090 ;
        RECT  1.870 2.265 1.965 3.205 ;
        END
        ANTENNADIFFAREA     0.7625 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 1.290 2.715 1.845 ;
        RECT  2.425 1.290 2.555 1.580 ;
        RECT  1.205 1.290 2.425 1.450 ;
        END
        ANTENNAGATEAREA     0.3185 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.540 0.480 2.000 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.635 1.310 2.035 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.005 -0.250 3.220 0.250 ;
        RECT  2.745 -0.250 3.005 0.745 ;
        RECT  1.265 -0.250 2.745 0.250 ;
        RECT  1.005 -0.250 1.265 0.860 ;
        RECT  0.000 -0.250 1.005 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.695 3.440 3.220 3.940 ;
        RECT  2.435 2.545 2.695 3.940 ;
        RECT  1.545 3.440 2.435 3.940 ;
        RECT  1.285 2.555 1.545 3.940 ;
        RECT  0.385 3.440 1.285 3.940 ;
        RECT  0.125 2.205 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.690 1.630 1.950 1.790 ;
        RECT  1.530 1.630 1.690 2.375 ;
        RECT  0.925 2.215 1.530 2.375 ;
        RECT  0.825 2.215 0.925 2.535 ;
        RECT  0.665 0.970 0.825 2.535 ;
        RECT  0.385 0.970 0.665 1.130 ;
        RECT  0.125 0.870 0.385 1.130 ;
    END
END OAI2BB1X2

MACRO OAI2BB1X1
    CLASS CORE ;
    FOREIGN OAI2BB1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.485 2.205 2.475 ;
        RECT  2.125 1.105 2.175 2.475 ;
        RECT  2.045 0.895 2.125 2.475 ;
        RECT  1.965 0.895 2.045 1.645 ;
        RECT  1.775 2.315 2.045 2.475 ;
        RECT  1.825 0.895 1.965 1.155 ;
        RECT  1.515 2.315 1.775 2.915 ;
        END
        ANTENNADIFFAREA     0.4433 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.290 1.435 1.665 ;
        END
        ANTENNAGATEAREA     0.1586 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.440 0.595 0.585 0.855 ;
        RECT  0.125 0.470 0.440 0.855 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.875 0.955 2.135 ;
        RECT  0.585 1.700 0.795 2.135 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 -0.250 2.300 0.250 ;
        RECT  1.005 -0.250 1.265 1.110 ;
        RECT  0.000 -0.250 1.005 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 3.440 2.300 3.940 ;
        RECT  1.575 3.285 2.175 3.940 ;
        RECT  1.235 3.440 1.575 3.940 ;
        RECT  0.975 2.895 1.235 3.940 ;
        RECT  0.385 3.440 0.975 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.705 1.850 1.865 2.135 ;
        RECT  1.335 1.975 1.705 2.135 ;
        RECT  1.175 1.975 1.335 2.475 ;
        RECT  0.785 2.315 1.175 2.475 ;
        RECT  0.525 2.315 0.785 2.575 ;
        RECT  0.385 2.315 0.525 2.475 ;
        RECT  0.225 1.035 0.385 2.475 ;
        RECT  0.125 1.035 0.225 1.295 ;
    END
END OAI2BB1X1

MACRO OAI2BB1XL
    CLASS CORE ;
    FOREIGN OAI2BB1XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 0.945 2.205 1.895 ;
        RECT  2.115 0.945 2.175 2.450 ;
        RECT  2.045 0.850 2.115 2.450 ;
        RECT  1.855 0.850 2.045 1.110 ;
        RECT  2.015 1.735 2.045 2.450 ;
        RECT  1.965 2.110 2.015 2.450 ;
        RECT  1.940 2.290 1.965 2.450 ;
        RECT  1.680 2.290 1.940 2.890 ;
        END
        ANTENNADIFFAREA     0.3867 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.985 1.290 1.375 1.615 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.440 0.595 0.585 0.855 ;
        RECT  0.125 0.470 0.440 0.855 ;
        END
        ANTENNAGATEAREA     0.0572 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.885 1.015 2.145 ;
        RECT  0.585 1.700 0.795 2.145 ;
        END
        ANTENNAGATEAREA     0.0572 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 -0.250 2.300 0.250 ;
        RECT  1.005 -0.250 1.265 1.110 ;
        RECT  0.000 -0.250 1.005 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.980 3.440 2.300 3.940 ;
        RECT  1.720 3.285 1.980 3.940 ;
        RECT  1.360 3.440 1.720 3.940 ;
        RECT  1.100 2.895 1.360 3.940 ;
        RECT  0.385 3.440 1.100 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.715 1.290 1.865 1.555 ;
        RECT  1.555 1.290 1.715 1.955 ;
        RECT  1.355 1.795 1.555 1.955 ;
        RECT  1.195 1.795 1.355 2.510 ;
        RECT  0.815 2.350 1.195 2.510 ;
        RECT  0.555 2.350 0.815 2.610 ;
        RECT  0.385 2.350 0.555 2.510 ;
        RECT  0.225 1.035 0.385 2.510 ;
        RECT  0.125 1.035 0.225 1.295 ;
    END
END OAI2BB1XL

MACRO OAI33X4
    CLASS CORE ;
    FOREIGN OAI33X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.305 0.970 1.465 2.570 ;
        RECT  1.205 0.970 1.305 1.130 ;
        RECT  1.205 1.700 1.305 2.570 ;
        RECT  1.045 1.700 1.205 2.400 ;
        END
        ANTENNADIFFAREA     0.7906 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.055 0.600 2.315 0.815 ;
        RECT  1.715 0.600 2.055 0.760 ;
        RECT  1.505 0.470 1.715 0.760 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.180 1.460 2.625 1.620 ;
        RECT  2.175 1.460 2.180 1.925 ;
        RECT  2.020 1.460 2.175 1.990 ;
        RECT  1.965 1.700 2.020 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.845 1.435 3.105 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.615 1.495 4.935 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.020 1.455 4.095 1.615 ;
        RECT  4.015 1.455 4.020 1.965 ;
        RECT  3.810 1.455 4.015 1.990 ;
        RECT  3.805 1.700 3.810 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.520 3.605 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 -0.250 5.060 0.250 ;
        RECT  2.625 -0.250 2.885 0.405 ;
        RECT  2.160 -0.250 2.625 0.250 ;
        RECT  1.900 -0.250 2.160 0.405 ;
        RECT  0.925 -0.250 1.900 0.250 ;
        RECT  0.665 -0.250 0.925 0.845 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.690 3.440 5.060 3.940 ;
        RECT  4.430 2.510 4.690 3.940 ;
        RECT  2.005 3.440 4.430 3.940 ;
        RECT  1.745 3.285 2.005 3.940 ;
        RECT  0.925 3.440 1.745 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.640 0.995 4.900 1.255 ;
        RECT  4.435 1.095 4.640 1.255 ;
        RECT  4.275 1.095 4.435 2.330 ;
        RECT  3.945 1.095 4.275 1.255 ;
        RECT  3.505 2.170 4.275 2.330 ;
        RECT  3.685 0.995 3.945 1.255 ;
        RECT  3.065 2.170 3.505 2.430 ;
        RECT  3.175 0.995 3.435 1.255 ;
        RECT  2.485 1.095 3.175 1.255 ;
        RECT  2.905 2.170 3.065 2.910 ;
        RECT  0.675 2.750 2.905 2.910 ;
        RECT  2.225 0.995 2.485 1.255 ;
        RECT  1.015 1.360 1.120 1.520 ;
        RECT  0.855 1.165 1.015 1.520 ;
        RECT  0.385 1.165 0.855 1.325 ;
        RECT  0.515 1.505 0.675 2.910 ;
        RECT  0.430 1.505 0.515 1.765 ;
        RECT  0.250 0.595 0.385 1.325 ;
        RECT  0.250 1.945 0.335 2.905 ;
        RECT  0.175 0.595 0.250 2.905 ;
        RECT  0.125 0.595 0.175 2.105 ;
        RECT  0.090 1.165 0.125 2.105 ;
    END
END OAI33X4

MACRO OAI33X2
    CLASS CORE ;
    FOREIGN OAI33X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.290 1.290 6.315 2.585 ;
        RECT  6.240 1.155 6.290 2.585 ;
        RECT  6.080 1.155 6.240 3.050 ;
        RECT  5.785 1.155 6.080 1.315 ;
        RECT  5.900 2.890 6.080 3.050 ;
        RECT  5.640 2.890 5.900 3.085 ;
        RECT  5.525 0.970 5.785 1.315 ;
        RECT  3.370 2.890 5.640 3.050 ;
        RECT  4.765 1.155 5.525 1.315 ;
        RECT  4.505 0.970 4.765 1.315 ;
        RECT  3.745 1.155 4.505 1.315 ;
        RECT  3.485 0.970 3.745 1.315 ;
        RECT  2.610 2.890 3.370 3.215 ;
        RECT  0.385 2.890 2.610 3.050 ;
        RECT  0.125 2.275 0.385 3.215 ;
        END
        ANTENNADIFFAREA     2.1773 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 1.430 1.745 2.030 ;
        END
        ANTENNAGATEAREA     0.4290 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 1.410 2.425 1.670 ;
        RECT  2.165 1.410 2.325 2.370 ;
        RECT  1.070 2.210 2.165 2.370 ;
        RECT  1.070 1.700 1.255 1.990 ;
        RECT  0.910 1.475 1.070 2.370 ;
        RECT  0.775 1.475 0.910 1.735 ;
        END
        ANTENNAGATEAREA     0.4316 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.665 1.765 2.910 2.075 ;
        RECT  2.650 1.765 2.665 2.710 ;
        RECT  2.505 1.915 2.650 2.710 ;
        RECT  0.725 2.550 2.505 2.710 ;
        RECT  0.565 1.930 0.725 2.710 ;
        RECT  0.550 1.930 0.565 2.090 ;
        RECT  0.470 1.580 0.550 2.090 ;
        RECT  0.390 1.355 0.470 2.090 ;
        RECT  0.335 1.355 0.390 1.840 ;
        RECT  0.290 1.290 0.335 1.840 ;
        RECT  0.125 1.290 0.290 1.580 ;
        END
        ANTENNAGATEAREA     0.4290 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.335 1.555 4.595 2.025 ;
        RECT  4.265 1.700 4.335 1.990 ;
        END
        ANTENNAGATEAREA     0.4186 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.095 1.495 5.420 1.655 ;
        RECT  4.935 1.495 5.095 2.370 ;
        RECT  3.865 2.210 4.935 2.370 ;
        RECT  3.915 1.700 4.015 1.990 ;
        RECT  3.865 1.495 3.915 1.990 ;
        RECT  3.705 1.495 3.865 2.370 ;
        RECT  3.655 1.495 3.705 1.655 ;
        END
        ANTENNAGATEAREA     0.4186 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.750 5.900 2.175 ;
        RECT  5.795 1.700 5.855 2.175 ;
        RECT  5.645 1.700 5.795 2.710 ;
        RECT  5.640 1.750 5.645 2.710 ;
        RECT  5.635 1.800 5.640 2.710 ;
        RECT  3.395 2.550 5.635 2.710 ;
        RECT  3.235 1.765 3.395 2.710 ;
        RECT  3.135 1.765 3.235 2.025 ;
        END
        ANTENNAGATEAREA     0.4186 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.835 -0.250 6.440 0.250 ;
        RECT  2.575 -0.250 2.835 0.405 ;
        RECT  1.735 -0.250 2.575 0.250 ;
        RECT  1.475 -0.250 1.735 0.405 ;
        RECT  0.785 -0.250 1.475 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 3.440 6.440 3.940 ;
        RECT  4.320 3.285 4.580 3.940 ;
        RECT  1.630 3.440 4.320 3.940 ;
        RECT  1.370 3.285 1.630 3.940 ;
        RECT  0.000 3.440 1.370 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.190 0.815 6.295 0.975 ;
        RECT  6.030 0.615 6.190 0.975 ;
        RECT  5.280 0.615 6.030 0.775 ;
        RECT  5.015 0.615 5.280 0.975 ;
        RECT  4.255 0.615 5.015 0.775 ;
        RECT  3.995 0.615 4.255 0.975 ;
        RECT  3.235 0.615 3.995 0.775 ;
        RECT  3.075 0.615 3.235 1.105 ;
        RECT  2.975 0.845 3.075 1.105 ;
        RECT  2.285 0.945 2.975 1.105 ;
        RECT  2.025 0.845 2.285 1.105 ;
        RECT  1.335 0.945 2.025 1.105 ;
        RECT  1.075 0.845 1.335 1.105 ;
        RECT  0.385 0.945 1.075 1.105 ;
        RECT  0.125 0.845 0.385 1.105 ;
    END
END OAI33X2

MACRO OAI33X1
    CLASS CORE ;
    FOREIGN OAI33X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 1.105 3.555 2.175 ;
        RECT  3.500 1.105 3.515 2.405 ;
        RECT  3.345 0.865 3.500 2.405 ;
        RECT  3.340 0.865 3.345 1.515 ;
        RECT  2.570 2.245 3.345 2.405 ;
        RECT  3.185 0.865 3.340 1.225 ;
        RECT  2.425 1.065 3.185 1.225 ;
        RECT  2.410 2.245 2.570 2.770 ;
        RECT  2.165 0.955 2.425 1.225 ;
        RECT  1.815 2.610 2.410 2.770 ;
        RECT  1.555 2.610 1.815 3.210 ;
        END
        ANTENNADIFFAREA     0.9898 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.330 0.515 1.720 ;
        RECT  0.125 1.290 0.335 1.720 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.965 1.465 1.065 1.725 ;
        RECT  0.805 1.465 0.965 2.270 ;
        RECT  0.795 2.110 0.805 2.270 ;
        RECT  0.585 2.110 0.795 2.400 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.350 1.790 1.575 2.170 ;
        RECT  1.315 1.790 1.350 2.745 ;
        RECT  1.255 2.010 1.315 2.745 ;
        RECT  1.190 2.010 1.255 2.810 ;
        RECT  1.045 2.520 1.190 2.810 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.845 1.585 3.105 2.055 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.460 2.635 1.990 ;
        RECT  2.345 1.460 2.425 1.880 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.055 2.110 2.175 2.400 ;
        RECT  1.895 1.465 2.055 2.400 ;
        RECT  1.795 1.465 1.895 1.725 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 -0.250 3.680 0.250 ;
        RECT  1.145 -0.250 1.405 0.935 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 0.940 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 3.440 3.680 3.940 ;
        RECT  2.760 2.835 3.020 3.940 ;
        RECT  0.470 3.440 2.760 3.940 ;
        RECT  0.210 2.615 0.470 3.940 ;
        RECT  0.000 3.440 0.210 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.675 0.615 2.935 0.885 ;
        RECT  1.915 0.615 2.675 0.775 ;
        RECT  1.815 0.615 1.915 1.125 ;
        RECT  1.755 0.615 1.815 1.280 ;
        RECT  1.655 0.865 1.755 1.280 ;
        RECT  0.895 1.120 1.655 1.280 ;
        RECT  0.735 0.845 0.895 1.280 ;
        RECT  0.635 0.845 0.735 1.105 ;
    END
END OAI33X1

MACRO OAI33XL
    CLASS CORE ;
    FOREIGN OAI33XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 0.880 3.555 2.175 ;
        RECT  3.505 0.880 3.515 2.330 ;
        RECT  3.345 0.740 3.505 2.330 ;
        RECT  3.245 0.740 3.345 1.270 ;
        RECT  1.755 2.170 3.345 2.330 ;
        RECT  2.515 1.110 3.245 1.270 ;
        RECT  2.355 0.810 2.515 1.270 ;
        RECT  2.195 0.810 2.355 0.970 ;
        RECT  1.495 2.170 1.755 2.430 ;
        END
        ANTENNADIFFAREA     0.5572 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.405 1.740 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.480 1.025 1.640 ;
        RECT  0.635 1.480 0.795 1.990 ;
        RECT  0.585 1.700 0.635 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.730 1.505 1.990 ;
        RECT  1.245 1.730 1.255 2.400 ;
        RECT  1.095 1.830 1.245 2.400 ;
        RECT  1.045 2.110 1.095 2.400 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.840 1.500 3.100 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.700 2.635 1.990 ;
        RECT  2.395 1.450 2.585 1.990 ;
        RECT  2.355 1.450 2.395 1.710 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.700 2.175 1.990 ;
        RECT  1.725 1.730 1.965 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 -0.250 3.680 0.250 ;
        RECT  1.145 -0.250 1.405 0.930 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.000 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.000 3.440 3.680 3.940 ;
        RECT  2.740 2.510 3.000 3.940 ;
        RECT  0.515 3.440 2.740 3.940 ;
        RECT  0.255 2.205 0.515 3.940 ;
        RECT  0.000 3.440 0.255 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.890 0.770 2.995 0.930 ;
        RECT  2.730 0.470 2.890 0.930 ;
        RECT  1.915 0.470 2.730 0.630 ;
        RECT  1.755 0.470 1.915 1.000 ;
        RECT  1.745 0.735 1.755 1.000 ;
        RECT  1.585 0.735 1.745 1.280 ;
        RECT  0.895 1.120 1.585 1.280 ;
        RECT  0.735 0.740 0.895 1.280 ;
        RECT  0.635 0.740 0.735 1.000 ;
    END
END OAI33XL

MACRO OAI32X4
    CLASS CORE ;
    FOREIGN OAI32X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.700 4.475 2.995 ;
        RECT  4.385 1.040 4.450 2.995 ;
        RECT  4.350 0.640 4.385 2.995 ;
        RECT  4.250 0.640 4.350 3.195 ;
        RECT  4.125 0.640 4.250 1.240 ;
        RECT  4.090 2.255 4.250 3.195 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 2.110 2.635 2.400 ;
        RECT  2.410 1.785 2.570 2.400 ;
        RECT  2.310 1.785 2.410 1.945 ;
        END
        ANTENNAGATEAREA     0.1092 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 2.520 2.175 2.810 ;
        RECT  1.965 2.520 2.150 2.935 ;
        RECT  1.715 2.675 1.965 2.935 ;
        END
        ANTENNAGATEAREA     0.1092 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.450 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.260 1.105 1.495 ;
        RECT  0.585 1.260 0.795 1.580 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 1.575 1.575 1.860 ;
        RECT  1.255 1.700 1.315 1.860 ;
        RECT  1.045 1.700 1.255 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.895 -0.250 5.060 0.250 ;
        RECT  4.635 -0.250 4.895 1.230 ;
        RECT  3.875 -0.250 4.635 0.250 ;
        RECT  3.615 -0.250 3.875 0.820 ;
        RECT  1.325 -0.250 3.615 0.250 ;
        RECT  1.065 -0.250 1.325 0.405 ;
        RECT  0.385 -0.250 1.065 0.250 ;
        RECT  0.125 -0.250 0.385 1.155 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.920 3.440 5.060 3.940 ;
        RECT  4.660 2.175 4.920 3.940 ;
        RECT  3.810 3.440 4.660 3.940 ;
        RECT  3.550 2.375 3.810 3.940 ;
        RECT  2.665 3.440 3.550 3.940 ;
        RECT  2.405 2.830 2.665 3.940 ;
        RECT  0.385 3.440 2.405 3.940 ;
        RECT  0.125 2.175 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.945 1.585 4.060 1.845 ;
        RECT  3.785 1.020 3.945 2.080 ;
        RECT  3.415 1.020 3.785 1.180 ;
        RECT  3.260 1.920 3.785 2.080 ;
        RECT  3.180 1.445 3.440 1.740 ;
        RECT  3.255 0.525 3.415 1.180 ;
        RECT  3.100 1.920 3.260 2.905 ;
        RECT  3.105 0.525 3.255 0.785 ;
        RECT  2.455 1.445 3.180 1.605 ;
        RECT  3.000 1.965 3.100 2.905 ;
        RECT  2.865 1.085 2.965 1.245 ;
        RECT  2.705 0.680 2.865 1.245 ;
        RECT  1.915 0.680 2.705 0.840 ;
        RECT  2.195 1.035 2.455 1.605 ;
        RECT  2.075 1.445 2.195 1.605 ;
        RECT  1.915 1.445 2.075 2.330 ;
        RECT  1.755 0.680 1.915 1.130 ;
        RECT  1.690 2.170 1.915 2.330 ;
        RECT  1.655 0.870 1.755 1.130 ;
        RECT  1.430 2.170 1.690 2.430 ;
        RECT  0.665 0.920 1.655 1.080 ;
    END
END OAI32X4

MACRO OAI32X2
    CLASS CORE ;
    FOREIGN OAI32X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.980 1.290 5.395 1.580 ;
        RECT  4.950 1.065 4.980 2.670 ;
        RECT  4.860 1.065 4.950 2.835 ;
        RECT  4.820 0.895 4.860 2.835 ;
        RECT  4.600 0.895 4.820 1.225 ;
        RECT  4.680 2.235 4.820 2.835 ;
        RECT  3.095 2.510 4.680 2.670 ;
        RECT  3.840 1.065 4.600 1.225 ;
        RECT  3.580 0.895 3.840 1.225 ;
        RECT  2.930 2.510 3.095 2.995 ;
        RECT  2.670 2.275 2.930 3.215 ;
        RECT  2.610 2.510 2.670 2.810 ;
        RECT  0.610 2.510 2.610 2.670 ;
        RECT  0.465 2.510 0.610 2.810 ;
        RECT  0.205 2.275 0.465 3.215 ;
        RECT  0.125 2.745 0.205 2.995 ;
        END
        ANTENNADIFFAREA     1.8920 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.885 1.530 4.130 1.990 ;
        RECT  3.805 1.700 3.885 1.990 ;
        END
        ANTENNAGATEAREA     0.3666 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.500 1.665 4.610 1.925 ;
        RECT  4.340 1.665 4.500 2.330 ;
        RECT  3.505 2.170 4.340 2.330 ;
        RECT  3.555 1.405 3.620 1.565 ;
        RECT  3.505 1.405 3.555 1.990 ;
        RECT  3.345 1.405 3.505 2.330 ;
        END
        ANTENNAGATEAREA     0.3666 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.500 1.680 1.715 1.990 ;
        RECT  1.245 1.760 1.500 1.990 ;
        END
        ANTENNAGATEAREA     0.4264 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 1.290 2.055 1.735 ;
        RECT  1.255 1.290 1.895 1.450 ;
        RECT  1.065 1.290 1.255 1.580 ;
        RECT  0.905 1.290 1.065 1.735 ;
        END
        ANTENNAGATEAREA     0.4316 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.430 1.790 2.990 2.050 ;
        RECT  2.270 1.790 2.430 2.330 ;
        RECT  0.950 2.170 2.270 2.330 ;
        RECT  0.790 1.930 0.950 2.330 ;
        RECT  0.635 1.930 0.790 2.090 ;
        RECT  0.475 1.395 0.635 2.090 ;
        RECT  0.335 1.395 0.475 1.655 ;
        RECT  0.125 1.290 0.335 1.655 ;
        END
        ANTENNAGATEAREA     0.4264 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.905 -0.250 5.520 0.250 ;
        RECT  2.645 -0.250 2.905 0.405 ;
        RECT  1.845 -0.250 2.645 0.250 ;
        RECT  1.585 -0.250 1.845 0.745 ;
        RECT  0.785 -0.250 1.585 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.980 3.440 5.520 3.940 ;
        RECT  3.720 2.895 3.980 3.940 ;
        RECT  1.645 3.440 3.720 3.940 ;
        RECT  1.385 2.895 1.645 3.940 ;
        RECT  0.000 3.440 1.385 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.110 0.555 5.370 0.885 ;
        RECT  4.350 0.555 5.110 0.715 ;
        RECT  4.090 0.555 4.350 0.885 ;
        RECT  3.330 0.555 4.090 0.715 ;
        RECT  3.170 0.555 3.330 1.085 ;
        RECT  3.070 0.790 3.170 1.085 ;
        RECT  2.355 0.925 3.070 1.085 ;
        RECT  2.095 0.685 2.355 1.085 ;
        RECT  1.335 0.925 2.095 1.085 ;
        RECT  1.175 0.675 1.335 1.085 ;
        RECT  1.075 0.675 1.175 0.935 ;
        RECT  0.385 0.775 1.075 0.935 ;
        RECT  0.125 0.775 0.385 1.035 ;
    END
END OAI32X2

MACRO OAI32X1
    CLASS CORE ;
    FOREIGN OAI32X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.515 1.515 2.635 1.990 ;
        RECT  2.355 0.895 2.515 2.330 ;
        RECT  2.255 0.895 2.355 1.155 ;
        RECT  1.715 2.170 2.355 2.330 ;
        RECT  1.695 2.170 1.715 2.585 ;
        RECT  1.435 2.040 1.695 2.980 ;
        END
        ANTENNADIFFAREA     0.8970 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.405 3.095 1.990 ;
        RECT  2.815 1.405 2.885 1.915 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.095 1.700 2.175 1.990 ;
        RECT  1.935 1.265 2.095 1.990 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.450 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.290 1.105 1.485 ;
        RECT  0.585 1.290 0.905 1.580 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.530 1.300 1.575 1.560 ;
        RECT  1.475 1.300 1.530 1.580 ;
        RECT  1.315 1.300 1.475 1.860 ;
        RECT  1.255 1.700 1.315 1.860 ;
        RECT  1.045 1.700 1.255 1.990 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 -0.250 3.220 0.250 ;
        RECT  1.205 -0.250 1.465 0.745 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 1.155 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.655 3.440 3.220 3.940 ;
        RECT  2.395 2.555 2.655 3.940 ;
        RECT  0.385 3.440 2.395 3.940 ;
        RECT  0.125 2.205 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.985 0.885 3.085 1.145 ;
        RECT  2.825 0.555 2.985 1.145 ;
        RECT  2.005 0.555 2.825 0.715 ;
        RECT  1.845 0.555 2.005 1.085 ;
        RECT  1.745 0.790 1.845 1.085 ;
        RECT  0.925 0.925 1.745 1.085 ;
        RECT  0.665 0.825 0.925 1.085 ;
    END
END OAI32X1

MACRO OAI32XL
    CLASS CORE ;
    FOREIGN OAI32XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.515 1.515 2.635 1.990 ;
        RECT  2.355 0.900 2.515 2.330 ;
        RECT  2.255 0.900 2.355 1.160 ;
        RECT  1.760 2.170 2.355 2.330 ;
        RECT  1.500 2.135 1.760 2.395 ;
        END
        ANTENNADIFFAREA     0.3742 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 1.480 3.095 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 1.700 2.175 1.990 ;
        RECT  1.965 1.345 2.145 1.990 ;
        RECT  1.885 1.345 1.965 1.505 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.470 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.290 1.105 1.515 ;
        RECT  0.585 1.290 0.905 1.580 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 1.300 1.575 1.560 ;
        RECT  1.315 1.300 1.475 1.860 ;
        RECT  1.255 1.700 1.315 1.860 ;
        RECT  1.045 1.700 1.255 1.990 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 -0.250 3.220 0.250 ;
        RECT  1.205 -0.250 1.465 0.750 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 1.170 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.655 3.440 3.220 3.940 ;
        RECT  2.395 2.555 2.655 3.940 ;
        RECT  0.540 3.440 2.395 3.940 ;
        RECT  0.280 2.175 0.540 3.940 ;
        RECT  0.000 3.440 0.280 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.035 1.030 3.085 1.290 ;
        RECT  2.875 0.555 3.035 1.290 ;
        RECT  2.005 0.555 2.875 0.715 ;
        RECT  2.825 1.030 2.875 1.290 ;
        RECT  1.845 0.555 2.005 1.110 ;
        RECT  0.665 0.950 1.845 1.110 ;
    END
END OAI32XL

MACRO OAI31X4
    CLASS CORE ;
    FOREIGN OAI31X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 1.290 4.475 1.990 ;
        RECT  4.225 1.095 4.465 2.295 ;
        RECT  4.015 1.095 4.225 1.335 ;
        RECT  3.805 2.055 4.225 2.295 ;
        RECT  3.955 0.695 4.015 1.335 ;
        RECT  3.695 0.595 3.955 1.335 ;
        RECT  3.545 2.055 3.805 3.065 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 2.110 2.255 2.585 ;
        END
        ANTENNAGATEAREA     0.0936 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.415 1.945 0.675 2.205 ;
        RECT  0.335 1.945 0.415 2.105 ;
        RECT  0.150 1.700 0.335 2.105 ;
        RECT  0.125 1.700 0.150 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.350 0.985 1.680 ;
        RECT  0.585 1.290 0.795 1.680 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.385 1.285 1.620 1.545 ;
        RECT  1.360 1.285 1.385 2.155 ;
        RECT  1.255 1.335 1.360 2.155 ;
        RECT  1.225 1.335 1.255 2.400 ;
        RECT  1.070 1.995 1.225 2.400 ;
        RECT  1.045 2.110 1.070 2.400 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 -0.250 4.600 0.250 ;
        RECT  4.205 -0.250 4.465 0.870 ;
        RECT  3.445 -0.250 4.205 0.250 ;
        RECT  3.185 -0.250 3.445 1.020 ;
        RECT  1.365 -0.250 3.185 0.250 ;
        RECT  1.105 -0.250 1.365 0.745 ;
        RECT  0.385 -0.250 1.105 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.315 3.440 4.600 3.940 ;
        RECT  4.055 2.505 4.315 3.940 ;
        RECT  3.295 3.440 4.055 3.940 ;
        RECT  3.035 2.480 3.295 3.940 ;
        RECT  2.275 3.440 3.035 3.940 ;
        RECT  2.015 2.850 2.275 3.940 ;
        RECT  0.505 3.440 2.015 3.940 ;
        RECT  0.245 2.550 0.505 3.940 ;
        RECT  0.000 3.440 0.245 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.355 1.555 3.690 1.815 ;
        RECT  3.195 1.240 3.355 2.275 ;
        RECT  2.935 1.240 3.195 1.400 ;
        RECT  2.785 2.115 3.195 2.275 ;
        RECT  2.675 0.695 2.935 1.400 ;
        RECT  2.370 1.635 2.930 1.895 ;
        RECT  2.525 2.115 2.785 3.085 ;
        RECT  2.370 0.860 2.425 1.120 ;
        RECT  2.210 0.860 2.370 1.895 ;
        RECT  2.165 0.860 2.210 1.120 ;
        RECT  1.755 1.735 2.210 1.895 ;
        RECT  1.655 0.840 1.915 1.100 ;
        RECT  1.595 1.735 1.755 2.900 ;
        RECT  0.815 0.940 1.655 1.100 ;
        RECT  1.395 2.640 1.595 2.900 ;
        RECT  0.555 0.840 0.815 1.100 ;
    END
END OAI31X4

MACRO OAI31X2
    CLASS CORE ;
    FOREIGN OAI31X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.995 1.515 4.015 2.515 ;
        RECT  3.805 0.955 3.995 2.515 ;
        RECT  3.695 0.955 3.805 1.215 ;
        RECT  3.655 2.355 3.805 2.515 ;
        RECT  3.495 2.355 3.655 2.865 ;
        RECT  3.395 2.605 3.495 2.865 ;
        RECT  1.925 2.605 3.395 2.765 ;
        RECT  1.665 2.585 1.925 3.185 ;
        END
        ANTENNADIFFAREA     0.8832 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.470 3.625 1.840 ;
        RECT  3.345 1.470 3.555 1.990 ;
        END
        ANTENNAGATEAREA     0.3172 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 1.625 3.145 2.395 ;
        RECT  2.885 1.625 3.095 2.400 ;
        RECT  1.280 2.235 2.885 2.395 ;
        RECT  1.120 1.865 1.280 2.395 ;
        RECT  1.045 1.865 1.120 2.175 ;
        RECT  0.750 1.865 1.045 2.025 ;
        RECT  0.490 1.770 0.750 2.030 ;
        END
        ANTENNAGATEAREA     0.4290 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.480 1.445 2.580 1.705 ;
        RECT  2.320 1.270 2.480 1.705 ;
        RECT  1.255 1.270 2.320 1.430 ;
        RECT  1.235 1.270 1.255 1.580 ;
        RECT  0.975 1.270 1.235 1.670 ;
        END
        ANTENNAGATEAREA     0.4290 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.675 1.965 1.990 ;
        RECT  1.505 1.700 1.540 1.990 ;
        END
        ANTENNAGATEAREA     0.4290 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 -0.250 4.600 0.250 ;
        RECT  2.675 -0.250 2.935 0.405 ;
        RECT  1.915 -0.250 2.675 0.250 ;
        RECT  1.655 -0.250 1.915 0.405 ;
        RECT  0.895 -0.250 1.655 0.250 ;
        RECT  0.635 -0.250 0.895 0.405 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.165 3.440 4.600 3.940 ;
        RECT  3.905 2.760 4.165 3.940 ;
        RECT  3.105 3.440 3.905 3.940 ;
        RECT  2.845 2.945 3.105 3.940 ;
        RECT  0.765 3.440 2.845 3.940 ;
        RECT  0.505 2.255 0.765 3.940 ;
        RECT  0.000 3.440 0.505 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.365 0.865 4.465 1.125 ;
        RECT  4.205 0.565 4.365 1.125 ;
        RECT  3.445 0.565 4.205 0.725 ;
        RECT  3.285 0.565 3.445 1.075 ;
        RECT  3.185 0.815 3.285 1.075 ;
        RECT  2.425 0.850 3.185 1.010 ;
        RECT  2.165 0.800 2.425 1.060 ;
        RECT  1.405 0.850 2.165 1.010 ;
        RECT  1.145 0.800 1.405 1.060 ;
        RECT  0.385 0.900 1.145 1.060 ;
        RECT  0.125 0.900 0.385 1.160 ;
    END
END OAI31X2

MACRO OAI31X1
    CLASS CORE ;
    FOREIGN OAI31X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 1.105 2.635 2.400 ;
        RECT  2.585 1.105 2.610 2.500 ;
        RECT  2.425 0.790 2.585 2.500 ;
        RECT  2.245 0.790 2.425 1.050 ;
        RECT  1.805 2.340 2.425 2.500 ;
        RECT  1.545 2.340 1.805 2.940 ;
        END
        ANTENNADIFFAREA     0.5439 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 1.290 2.175 1.765 ;
        RECT  1.885 1.285 2.145 1.920 ;
        END
        ANTENNAGATEAREA     0.1586 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.790 0.675 2.050 ;
        RECT  0.125 1.700 0.335 2.050 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 1.420 1.155 1.710 ;
        RECT  0.795 1.420 0.895 1.580 ;
        RECT  0.585 1.290 0.795 1.580 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.535 1.635 1.635 1.895 ;
        RECT  1.375 1.635 1.535 2.115 ;
        RECT  1.255 1.955 1.375 2.115 ;
        RECT  1.070 1.955 1.255 2.400 ;
        RECT  1.045 2.110 1.070 2.400 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 -0.250 2.760 0.250 ;
        RECT  1.185 -0.250 1.445 0.405 ;
        RECT  0.385 -0.250 1.185 0.250 ;
        RECT  0.125 -0.250 0.385 1.155 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.315 3.440 2.760 3.940 ;
        RECT  2.055 2.680 2.315 3.940 ;
        RECT  0.675 3.440 2.055 3.940 ;
        RECT  0.415 2.270 0.675 3.940 ;
        RECT  0.000 3.440 0.415 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.735 0.820 1.995 1.080 ;
        RECT  0.895 0.870 1.735 1.030 ;
        RECT  0.635 0.770 0.895 1.030 ;
    END
END OAI31X1

MACRO OAI31XL
    CLASS CORE ;
    FOREIGN OAI31XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.015 0.490 2.175 2.810 ;
        RECT  1.965 0.490 2.015 1.355 ;
        RECT  1.965 2.520 2.015 2.810 ;
        RECT  1.915 0.490 1.965 0.650 ;
        RECT  1.625 2.635 1.965 2.795 ;
        RECT  1.365 2.635 1.625 2.895 ;
        END
        ANTENNADIFFAREA     0.4360 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.695 1.800 2.210 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 2.035 0.515 2.295 ;
        RECT  0.335 1.845 0.465 2.295 ;
        RECT  0.125 1.700 0.335 2.295 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.940 1.720 1.040 1.980 ;
        RECT  0.795 1.720 0.940 2.680 ;
        RECT  0.780 1.720 0.795 2.810 ;
        RECT  0.585 2.520 0.780 2.810 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 0.530 1.565 0.790 ;
        RECT  1.045 0.470 1.255 0.790 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.250 2.300 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 3.440 2.300 3.940 ;
        RECT  1.915 3.285 2.175 3.940 ;
        RECT  0.385 3.440 1.915 3.940 ;
        RECT  0.125 2.625 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.475 1.035 1.735 1.295 ;
        RECT  0.785 1.085 1.475 1.245 ;
        RECT  0.575 0.845 0.785 1.245 ;
        RECT  0.525 0.845 0.575 1.105 ;
    END
END OAI31XL

MACRO OAI222X4
    CLASS CORE ;
    FOREIGN OAI222X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.290 1.290 5.395 1.990 ;
        RECT  5.050 1.290 5.290 2.310 ;
        RECT  4.935 1.290 5.050 1.530 ;
        RECT  4.935 2.070 5.050 2.310 ;
        RECT  4.885 0.695 4.935 1.530 ;
        RECT  4.885 2.070 4.935 2.995 ;
        RECT  4.645 0.530 4.885 1.530 ;
        RECT  4.625 2.070 4.885 3.110 ;
        RECT  4.625 0.530 4.645 1.230 ;
        END
        ANTENNADIFFAREA     0.7688 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.505 2.650 1.975 ;
        RECT  2.425 1.505 2.635 1.990 ;
        RECT  2.390 1.505 2.425 1.975 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.390 1.615 3.635 1.990 ;
        RECT  3.230 1.615 3.390 2.090 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.460 2.195 0.720 2.455 ;
        RECT  0.365 2.195 0.460 2.400 ;
        RECT  0.335 1.765 0.365 2.400 ;
        RECT  0.310 1.700 0.335 2.400 ;
        RECT  0.205 1.700 0.310 2.355 ;
        RECT  0.125 1.700 0.205 2.175 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.715 1.170 1.990 ;
        RECT  0.585 1.700 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 2.200 2.360 2.520 ;
        RECT  1.965 2.110 2.175 2.520 ;
        RECT  1.935 2.200 1.965 2.520 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.460 1.750 1.935 ;
        RECT  1.505 1.460 1.715 1.990 ;
        RECT  1.405 1.460 1.505 1.935 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 -0.250 5.520 0.250 ;
        RECT  5.135 -0.250 5.395 1.080 ;
        RECT  4.335 -0.250 5.135 0.250 ;
        RECT  4.075 -0.250 4.335 0.405 ;
        RECT  1.100 -0.250 4.075 0.250 ;
        RECT  0.840 -0.250 1.100 0.405 ;
        RECT  0.805 1.230 1.065 1.520 ;
        RECT  0.500 -0.250 0.840 0.250 ;
        RECT  0.500 1.230 0.805 1.490 ;
        RECT  0.240 -0.250 0.500 1.490 ;
        RECT  0.000 -0.250 0.240 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 3.440 5.520 3.940 ;
        RECT  5.135 2.560 5.395 3.940 ;
        RECT  4.375 3.440 5.135 3.940 ;
        RECT  4.115 2.570 4.375 3.940 ;
        RECT  2.415 3.440 4.115 3.940 ;
        RECT  2.155 3.285 2.415 3.940 ;
        RECT  0.720 3.440 2.155 3.940 ;
        RECT  0.460 2.700 0.720 3.940 ;
        RECT  0.000 3.440 0.460 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.405 1.725 4.775 1.885 ;
        RECT  4.245 0.920 4.405 2.380 ;
        RECT  3.940 0.920 4.245 1.080 ;
        RECT  3.865 2.220 4.245 2.380 ;
        RECT  3.900 1.260 4.060 1.895 ;
        RECT  3.680 0.820 3.940 1.080 ;
        RECT  3.030 1.260 3.900 1.420 ;
        RECT  3.605 2.220 3.865 3.180 ;
        RECT  3.020 2.575 3.275 2.920 ;
        RECT  3.020 0.985 3.030 1.420 ;
        RECT  2.860 0.985 3.020 2.920 ;
        RECT  2.770 0.985 2.860 1.245 ;
        RECT  1.540 2.760 2.860 2.920 ;
        RECT  1.990 0.970 2.080 1.230 ;
        RECT  1.820 0.845 1.990 1.230 ;
        RECT  1.040 0.845 1.820 1.005 ;
        RECT  1.280 2.660 1.540 2.920 ;
        RECT  0.780 0.745 1.040 1.005 ;
    END
END OAI222X4

MACRO OAI222X2
    CLASS CORE ;
    FOREIGN OAI222X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.630 1.515 6.775 2.585 ;
        RECT  6.470 1.280 6.630 2.745 ;
        RECT  6.185 1.280 6.470 1.585 ;
        RECT  5.425 2.585 6.470 2.745 ;
        RECT  5.950 1.020 6.185 1.585 ;
        RECT  5.925 1.020 5.950 1.315 ;
        RECT  5.165 1.155 5.925 1.315 ;
        RECT  5.165 2.585 5.425 2.910 ;
        RECT  4.905 1.020 5.165 1.315 ;
        RECT  3.835 2.585 5.165 2.745 ;
        RECT  3.405 2.585 3.835 2.910 ;
        RECT  1.990 2.585 3.405 2.745 ;
        RECT  1.615 2.585 1.990 2.845 ;
        END
        ANTENNADIFFAREA     1.4676 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.135 1.930 6.245 2.190 ;
        RECT  5.975 1.930 6.135 2.405 ;
        RECT  4.935 2.245 5.975 2.405 ;
        RECT  4.885 1.925 4.935 2.405 ;
        RECT  4.725 1.655 4.885 2.405 ;
        RECT  4.600 1.655 4.725 1.915 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 1.590 5.650 1.990 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.430 1.665 2.530 1.925 ;
        RECT  2.270 1.665 2.430 2.395 ;
        RECT  1.585 2.235 2.270 2.395 ;
        RECT  1.425 2.140 1.585 2.395 ;
        RECT  0.795 2.140 1.425 2.300 ;
        RECT  0.755 1.685 0.795 2.300 ;
        RECT  0.635 1.635 0.755 2.300 ;
        RECT  0.585 1.635 0.635 1.990 ;
        RECT  0.495 1.635 0.585 1.895 ;
        END
        ANTENNAGATEAREA     0.3744 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 1.795 2.050 2.055 ;
        RECT  1.220 1.795 1.790 1.955 ;
        RECT  1.220 1.290 1.255 1.580 ;
        RECT  1.060 1.290 1.220 1.955 ;
        RECT  1.045 1.290 1.060 1.580 ;
        END
        ANTENNAGATEAREA     0.3744 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.070 1.905 4.315 2.165 ;
        RECT  3.910 1.905 4.070 2.405 ;
        RECT  3.805 2.110 3.910 2.405 ;
        RECT  3.010 2.245 3.805 2.405 ;
        RECT  2.850 1.720 3.010 2.405 ;
        RECT  2.750 1.720 2.850 1.980 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.565 3.620 2.050 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.285 -0.250 6.900 0.250 ;
        RECT  2.025 -0.250 2.285 0.405 ;
        RECT  1.450 -0.250 2.025 0.250 ;
        RECT  1.190 -0.250 1.450 0.405 ;
        RECT  0.390 -0.250 1.190 0.250 ;
        RECT  0.130 -0.250 0.390 1.015 ;
        RECT  0.000 -0.250 0.130 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.285 3.440 6.900 3.940 ;
        RECT  6.025 2.945 6.285 3.940 ;
        RECT  4.545 3.440 6.025 3.940 ;
        RECT  4.285 2.935 4.545 3.940 ;
        RECT  2.765 3.440 4.285 3.940 ;
        RECT  2.505 2.945 2.765 3.940 ;
        RECT  1.015 3.440 2.505 3.940 ;
        RECT  0.755 2.525 1.015 3.940 ;
        RECT  0.000 3.440 0.755 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.435 0.630 6.695 1.050 ;
        RECT  5.675 0.630 6.435 0.790 ;
        RECT  5.415 0.630 5.675 0.945 ;
        RECT  4.655 0.630 5.415 0.790 ;
        RECT  4.495 0.630 4.655 1.250 ;
        RECT  4.395 0.990 4.495 1.250 ;
        RECT  3.885 0.940 4.145 1.540 ;
        RECT  3.145 1.160 3.885 1.320 ;
        RECT  2.985 0.940 3.145 1.540 ;
        RECT  1.885 1.160 2.985 1.320 ;
        RECT  1.725 0.830 1.885 1.320 ;
        RECT  1.625 0.830 1.725 1.090 ;
        RECT  0.900 0.830 1.625 0.990 ;
        RECT  0.640 0.775 0.900 1.035 ;
    END
END OAI222X2

MACRO OAI222X1
    CLASS CORE ;
    FOREIGN OAI222X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.995 1.290 4.015 2.570 ;
        RECT  3.855 1.130 3.995 2.570 ;
        RECT  3.805 1.130 3.855 1.580 ;
        RECT  3.830 2.335 3.855 2.570 ;
        RECT  3.615 2.410 3.830 2.570 ;
        RECT  3.485 1.130 3.805 1.290 ;
        RECT  3.355 2.410 3.615 3.010 ;
        RECT  3.225 1.030 3.485 1.290 ;
        RECT  3.345 2.745 3.355 3.010 ;
        RECT  1.910 2.850 3.345 3.010 ;
        RECT  1.650 2.750 1.910 3.010 ;
        END
        ANTENNADIFFAREA     0.8640 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 1.485 3.135 1.745 ;
        RECT  2.885 1.485 3.095 2.400 ;
        RECT  2.875 1.485 2.885 1.765 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.735 3.645 2.150 ;
        RECT  3.345 1.700 3.555 2.150 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.350 2.170 0.600 2.430 ;
        RECT  0.125 1.970 0.350 2.430 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.470 1.065 1.730 ;
        RECT  0.585 1.470 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.305 1.820 2.565 2.270 ;
        RECT  2.175 2.110 2.305 2.270 ;
        RECT  1.965 2.110 2.175 2.400 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.470 2.085 1.730 ;
        RECT  1.505 1.470 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 -0.250 4.140 0.250 ;
        RECT  1.185 -0.250 1.445 0.865 ;
        RECT  0.385 -0.250 1.185 0.250 ;
        RECT  0.125 -0.250 0.385 1.275 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.765 3.440 4.140 3.940 ;
        RECT  2.505 3.285 2.765 3.940 ;
        RECT  1.040 3.440 2.505 3.940 ;
        RECT  0.780 2.430 1.040 3.940 ;
        RECT  0.000 3.440 0.780 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.735 0.680 3.995 0.940 ;
        RECT  2.975 0.680 3.735 0.840 ;
        RECT  2.715 0.680 2.975 1.280 ;
        RECT  1.955 0.680 2.715 0.840 ;
        RECT  2.205 1.025 2.465 1.285 ;
        RECT  0.895 1.125 2.205 1.285 ;
        RECT  1.695 0.680 1.955 0.940 ;
        RECT  0.635 0.675 0.895 1.285 ;
    END
END OAI222X1

MACRO OAI222XL
    CLASS CORE ;
    FOREIGN OAI222XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 1.290 3.555 2.585 ;
        RECT  3.275 1.075 3.435 2.875 ;
        RECT  3.155 1.075 3.275 1.235 ;
        RECT  2.970 2.615 3.275 2.875 ;
        RECT  2.895 0.975 3.155 1.235 ;
        RECT  1.530 2.715 2.970 2.875 ;
        RECT  1.245 2.580 1.530 2.875 ;
        END
        ANTENNADIFFAREA     0.4680 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.415 2.880 1.675 ;
        RECT  2.425 1.290 2.635 1.675 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.800 1.855 3.095 2.400 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.470 0.525 1.835 ;
        RECT  0.125 1.470 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.865 1.415 1.035 1.675 ;
        RECT  0.795 1.415 0.865 2.270 ;
        RECT  0.705 1.415 0.795 2.400 ;
        RECT  0.585 2.110 0.705 2.400 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.155 2.110 2.175 2.400 ;
        RECT  1.895 2.025 2.155 2.400 ;
        RECT  1.755 2.140 1.895 2.400 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.585 1.525 1.845 1.785 ;
        RECT  1.495 1.625 1.585 1.785 ;
        RECT  1.335 1.625 1.495 2.270 ;
        RECT  1.255 2.110 1.335 2.270 ;
        RECT  1.045 2.110 1.255 2.400 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.295 -0.250 3.680 0.250 ;
        RECT  1.035 -0.250 1.295 0.405 ;
        RECT  0.385 -0.250 1.035 0.250 ;
        RECT  0.125 -0.250 0.385 1.255 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.365 3.440 3.680 3.940 ;
        RECT  2.105 3.285 2.365 3.940 ;
        RECT  0.645 3.440 2.105 3.940 ;
        RECT  0.385 2.685 0.645 3.940 ;
        RECT  0.000 3.440 0.385 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.945 1.035 2.205 1.295 ;
        RECT  0.895 1.035 1.945 1.195 ;
        RECT  0.635 0.975 0.895 1.235 ;
    END
END OAI222XL

MACRO OAI221X4
    CLASS CORE ;
    FOREIGN OAI221X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 1.515 4.935 2.400 ;
        RECT  4.725 1.260 4.885 2.400 ;
        RECT  4.475 1.260 4.725 1.420 ;
        RECT  4.475 2.115 4.725 2.400 ;
        RECT  4.425 0.695 4.475 1.420 ;
        RECT  4.425 2.115 4.475 2.585 ;
        RECT  4.265 0.480 4.425 1.420 ;
        RECT  4.165 2.115 4.425 3.055 ;
        RECT  4.165 0.480 4.265 1.080 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.840 2.745 2.060 ;
        RECT  2.625 1.700 2.635 2.060 ;
        RECT  2.385 1.520 2.625 2.060 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.420 0.445 1.680 ;
        RECT  0.335 1.420 0.345 1.925 ;
        RECT  0.185 1.420 0.335 1.990 ;
        RECT  0.125 1.700 0.185 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.635 0.995 1.895 ;
        RECT  0.635 1.635 0.795 2.400 ;
        RECT  0.585 2.110 0.635 2.400 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 2.110 2.175 2.400 ;
        RECT  1.965 1.840 2.045 2.400 ;
        RECT  1.785 1.840 1.965 2.335 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 1.760 1.505 2.020 ;
        RECT  1.255 1.760 1.405 2.335 ;
        RECT  1.245 1.760 1.255 2.400 ;
        RECT  1.045 2.110 1.245 2.400 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 -0.250 5.060 0.250 ;
        RECT  4.675 -0.250 4.935 1.075 ;
        RECT  3.865 -0.250 4.675 0.250 ;
        RECT  3.705 -0.250 3.865 1.075 ;
        RECT  1.185 -0.250 3.705 0.250 ;
        RECT  0.925 -0.250 1.185 0.405 ;
        RECT  0.385 -0.250 0.925 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 3.440 5.060 3.940 ;
        RECT  4.675 2.595 4.935 3.940 ;
        RECT  3.865 3.440 4.675 3.940 ;
        RECT  3.705 2.565 3.865 3.940 ;
        RECT  3.590 3.285 3.705 3.940 ;
        RECT  3.005 3.440 3.590 3.940 ;
        RECT  2.745 3.285 3.005 3.940 ;
        RECT  1.945 3.440 2.745 3.940 ;
        RECT  1.685 3.285 1.945 3.940 ;
        RECT  0.385 3.440 1.685 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.525 1.630 4.420 1.790 ;
        RECT  3.405 0.915 3.525 2.845 ;
        RECT  3.365 0.475 3.405 2.845 ;
        RECT  3.145 0.475 3.365 1.075 ;
        RECT  3.145 2.685 3.365 2.845 ;
        RECT  3.020 1.475 3.180 2.485 ;
        RECT  2.995 1.475 3.020 1.635 ;
        RECT  2.545 2.325 3.020 2.485 ;
        RECT  2.835 1.375 2.995 1.635 ;
        RECT  2.385 2.325 2.545 3.130 ;
        RECT  2.235 2.705 2.385 3.130 ;
        RECT  1.165 2.705 2.235 2.865 ;
        RECT  1.995 1.280 2.095 1.540 ;
        RECT  1.835 1.035 1.995 1.540 ;
        RECT  0.785 1.035 1.835 1.195 ;
        RECT  0.905 2.605 1.165 2.865 ;
        RECT  0.525 0.985 0.785 1.245 ;
    END
END OAI221X4

MACRO OAI221X2
    CLASS CORE ;
    FOREIGN OAI221X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.895 2.110 4.935 2.400 ;
        RECT  4.735 1.290 4.895 2.560 ;
        RECT  4.425 1.290 4.735 1.450 ;
        RECT  4.725 2.110 4.735 2.560 ;
        RECT  4.385 2.400 4.725 2.560 ;
        RECT  4.265 1.030 4.425 1.450 ;
        RECT  4.125 2.400 4.385 2.900 ;
        RECT  4.165 1.030 4.265 1.290 ;
        RECT  3.435 2.400 4.125 2.560 ;
        RECT  3.275 2.400 3.435 2.775 ;
        RECT  3.095 2.615 3.275 2.775 ;
        RECT  2.940 2.615 3.095 2.995 ;
        RECT  2.680 2.615 2.940 3.215 ;
        RECT  1.300 2.615 2.680 2.775 ;
        RECT  1.040 2.585 1.300 2.845 ;
        END
        ANTENNADIFFAREA     1.1656 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.700 4.555 1.960 ;
        RECT  4.265 1.700 4.475 1.990 ;
        RECT  3.955 1.700 4.265 1.960 ;
        END
        ANTENNAGATEAREA     0.3380 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 1.610 2.055 1.770 ;
        RECT  1.680 1.610 1.840 2.360 ;
        RECT  0.610 2.200 1.680 2.360 ;
        RECT  0.545 2.175 0.610 2.360 ;
        RECT  0.385 1.635 0.545 2.360 ;
        RECT  0.285 1.635 0.385 1.990 ;
        RECT  0.125 1.700 0.285 1.990 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.855 1.635 1.385 1.990 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.960 3.590 2.220 ;
        RECT  3.330 1.685 3.555 2.220 ;
        RECT  2.400 1.685 3.330 1.845 ;
        RECT  2.290 1.685 2.400 2.205 ;
        RECT  2.240 1.685 2.290 2.305 ;
        RECT  2.030 2.045 2.240 2.305 ;
        END
        ANTENNAGATEAREA     0.3887 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 2.085 3.095 2.400 ;
        RECT  2.630 2.035 2.890 2.400 ;
        END
        ANTENNAGATEAREA     0.3887 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.465 -0.250 5.060 0.250 ;
        RECT  2.205 -0.250 2.465 0.405 ;
        RECT  1.405 -0.250 2.205 0.250 ;
        RECT  1.145 -0.250 1.405 1.030 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.290 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.895 3.440 5.060 3.940 ;
        RECT  4.635 2.755 4.895 3.940 ;
        RECT  3.875 3.440 4.635 3.940 ;
        RECT  3.615 2.755 3.875 3.940 ;
        RECT  2.120 3.440 3.615 3.940 ;
        RECT  1.860 2.955 2.120 3.940 ;
        RECT  0.385 3.440 1.860 3.940 ;
        RECT  0.125 2.640 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.835 0.800 4.935 1.060 ;
        RECT  4.675 0.655 4.835 1.060 ;
        RECT  3.915 0.655 4.675 0.815 ;
        RECT  3.655 0.520 3.915 1.290 ;
        RECT  2.895 0.520 3.655 0.680 ;
        RECT  3.145 0.890 3.405 1.490 ;
        RECT  1.915 1.240 3.145 1.400 ;
        RECT  2.735 0.520 2.895 1.010 ;
        RECT  2.635 0.750 2.735 1.010 ;
        RECT  1.655 0.690 1.915 1.400 ;
        RECT  0.895 1.240 1.655 1.400 ;
        RECT  0.635 0.690 0.895 1.400 ;
    END
END OAI221X2

MACRO OAI221X1
    CLASS CORE ;
    FOREIGN OAI221X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.490 1.105 3.555 2.400 ;
        RECT  3.330 0.665 3.490 2.400 ;
        RECT  3.230 0.665 3.330 1.265 ;
        RECT  3.095 2.215 3.330 2.400 ;
        RECT  3.090 2.215 3.095 2.585 ;
        RECT  2.830 2.215 3.090 2.895 ;
        RECT  1.715 2.215 2.830 2.375 ;
        RECT  1.595 2.215 1.715 2.995 ;
        RECT  1.435 2.215 1.595 3.190 ;
        RECT  1.335 2.590 1.435 3.190 ;
        END
        ANTENNADIFFAREA     0.7646 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.545 3.150 2.035 ;
        END
        ANTENNAGATEAREA     0.1703 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.720 0.495 2.130 ;
        RECT  0.125 1.700 0.335 2.130 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.205 1.925 1.255 2.400 ;
        RECT  1.085 1.735 1.205 2.400 ;
        RECT  1.045 1.635 1.085 2.400 ;
        RECT  0.825 1.635 1.045 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.350 1.475 2.635 2.020 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.475 1.785 2.035 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 -0.250 3.680 0.250 ;
        RECT  1.185 -0.250 1.445 0.405 ;
        RECT  0.385 -0.250 1.185 0.250 ;
        RECT  0.125 -0.250 0.385 1.290 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 3.440 3.680 3.940 ;
        RECT  2.225 2.555 2.485 3.940 ;
        RECT  0.735 3.440 2.225 3.940 ;
        RECT  0.475 2.500 0.735 3.940 ;
        RECT  0.000 3.440 0.475 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.720 0.695 2.980 1.295 ;
        RECT  1.960 1.135 2.720 1.295 ;
        RECT  2.210 0.660 2.470 0.955 ;
        RECT  0.895 0.660 2.210 0.820 ;
        RECT  1.700 1.035 1.960 1.295 ;
        RECT  0.635 0.660 0.895 1.260 ;
    END
END OAI221X1

MACRO OAI221XL
    CLASS CORE ;
    FOREIGN OAI221XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 1.105 3.095 2.810 ;
        RECT  3.045 1.030 3.080 2.810 ;
        RECT  2.910 1.030 3.045 2.910 ;
        RECT  2.885 1.030 2.910 2.960 ;
        RECT  2.820 1.030 2.885 1.290 ;
        RECT  2.590 2.700 2.885 2.960 ;
        RECT  1.530 2.740 2.590 2.900 ;
        RECT  1.195 2.695 1.530 2.955 ;
        END
        ANTENNADIFFAREA     0.4128 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 2.245 2.680 2.520 ;
        RECT  2.425 2.110 2.635 2.520 ;
        RECT  2.195 2.245 2.425 2.520 ;
        END
        ANTENNAGATEAREA     0.0910 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.220 0.480 2.530 ;
        RECT  0.125 2.110 0.335 2.530 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.685 1.350 1.895 ;
        RECT  0.585 1.685 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.495 2.400 1.755 ;
        RECT  1.965 1.495 2.175 1.990 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 2.110 1.650 2.395 ;
        RECT  1.045 2.110 1.255 2.400 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.010 -0.250 3.220 0.250 ;
        RECT  0.475 1.185 1.045 1.445 ;
        RECT  0.750 -0.250 1.010 0.405 ;
        RECT  0.475 -0.250 0.750 0.250 ;
        RECT  0.215 -0.250 0.475 1.445 ;
        RECT  0.000 -0.250 0.215 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.310 3.440 3.220 3.940 ;
        RECT  2.050 3.285 2.310 3.940 ;
        RECT  0.595 3.440 2.050 3.940 ;
        RECT  0.335 2.825 0.595 3.940 ;
        RECT  0.000 3.440 0.335 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.310 1.020 2.570 1.280 ;
        RECT  1.620 1.120 2.310 1.280 ;
        RECT  1.460 1.120 1.620 1.505 ;
        RECT  1.360 1.245 1.460 1.505 ;
    END
END OAI221XL

MACRO OAI22X4
    CLASS CORE ;
    FOREIGN OAI22X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.255 1.515 6.315 2.175 ;
        RECT  6.055 1.005 6.255 2.310 ;
        RECT  3.485 1.005 6.055 1.205 ;
        RECT  5.855 2.110 6.055 2.310 ;
        RECT  5.645 2.110 5.855 2.810 ;
        RECT  5.520 2.180 5.645 2.780 ;
        RECT  4.080 2.580 5.520 2.780 ;
        RECT  3.820 2.580 4.080 3.215 ;
        RECT  3.805 2.580 3.820 2.995 ;
        RECT  3.535 2.580 3.805 2.780 ;
        RECT  3.335 2.275 3.535 2.780 ;
        RECT  2.240 2.275 3.335 2.475 ;
        RECT  1.980 2.275 2.240 3.215 ;
        RECT  1.965 2.580 1.980 2.995 ;
        RECT  0.610 2.580 1.965 2.780 ;
        RECT  0.585 2.520 0.610 2.780 ;
        RECT  0.525 2.520 0.585 3.215 ;
        RECT  0.265 2.275 0.525 3.215 ;
        RECT  0.125 2.745 0.265 2.995 ;
        END
        ANTENNADIFFAREA     2.4653 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.690 1.615 2.950 1.875 ;
        RECT  2.675 1.615 2.690 1.775 ;
        RECT  2.515 1.495 2.675 1.775 ;
        RECT  1.305 1.495 2.515 1.655 ;
        RECT  1.255 1.495 1.305 1.825 ;
        RECT  1.045 1.495 1.255 1.990 ;
        END
        ANTENNAGATEAREA     0.7098 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.835 2.065 1.995 ;
        RECT  1.555 1.835 1.715 2.400 ;
        RECT  1.505 2.110 1.555 2.400 ;
        RECT  0.865 2.170 1.505 2.330 ;
        RECT  0.705 1.880 0.865 2.330 ;
        RECT  0.610 1.880 0.705 2.040 ;
        RECT  0.345 1.775 0.610 2.040 ;
        RECT  0.295 1.775 0.345 2.035 ;
        END
        ANTENNAGATEAREA     0.7098 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.870 1.825 5.130 2.400 ;
        RECT  4.725 2.110 4.870 2.400 ;
        RECT  3.875 2.240 4.725 2.400 ;
        RECT  3.715 1.730 3.875 2.400 ;
        RECT  3.530 1.730 3.715 1.990 ;
        RECT  3.430 1.730 3.530 1.890 ;
        RECT  3.170 1.630 3.430 1.890 ;
        END
        ANTENNAGATEAREA     0.7098 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.715 1.465 5.875 1.815 ;
        RECT  4.475 1.465 5.715 1.625 ;
        RECT  4.265 1.465 4.475 1.990 ;
        RECT  4.055 1.465 4.265 1.725 ;
        END
        ANTENNAGATEAREA     0.7098 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.685 -0.250 6.440 0.250 ;
        RECT  2.425 -0.250 2.685 0.405 ;
        RECT  1.885 -0.250 2.425 0.250 ;
        RECT  1.625 -0.250 1.885 0.405 ;
        RECT  0.935 -0.250 1.625 0.250 ;
        RECT  0.675 -0.250 0.935 0.405 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.930 3.440 6.440 3.940 ;
        RECT  4.670 2.960 4.930 3.940 ;
        RECT  3.150 3.440 4.670 3.940 ;
        RECT  2.890 2.655 3.150 3.940 ;
        RECT  1.380 3.440 2.890 3.940 ;
        RECT  1.120 2.960 1.380 3.940 ;
        RECT  0.000 3.440 1.120 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.235 0.665 6.295 0.825 ;
        RECT  2.975 0.665 3.235 1.375 ;
        RECT  2.285 1.155 2.975 1.315 ;
        RECT  2.025 1.055 2.285 1.315 ;
        RECT  1.335 1.155 2.025 1.315 ;
        RECT  1.075 1.025 1.335 1.315 ;
        RECT  0.385 1.155 1.075 1.315 ;
        RECT  0.125 0.695 0.385 1.315 ;
    END
END OAI22X4

MACRO OAI22X2
    CLASS CORE ;
    FOREIGN OAI22X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.425 1.515 4.475 2.585 ;
        RECT  4.265 1.200 4.425 2.700 ;
        RECT  3.955 1.200 4.265 1.360 ;
        RECT  2.935 2.540 4.265 2.700 ;
        RECT  3.695 0.955 3.955 1.360 ;
        RECT  2.935 1.200 3.695 1.360 ;
        RECT  2.775 0.955 2.935 1.360 ;
        RECT  2.610 2.540 2.935 2.965 ;
        RECT  2.675 0.955 2.775 1.215 ;
        RECT  1.235 2.540 2.610 2.700 ;
        RECT  1.075 2.540 1.235 2.965 ;
        RECT  0.975 2.705 1.075 2.965 ;
        END
        ANTENNADIFFAREA     1.0716 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 1.665 1.885 1.925 ;
        RECT  1.625 1.665 1.785 2.360 ;
        RECT  0.370 2.200 1.625 2.360 ;
        RECT  0.335 1.705 0.370 2.360 ;
        RECT  0.210 1.700 0.335 2.360 ;
        RECT  0.125 1.700 0.210 2.175 ;
        RECT  0.110 1.705 0.125 1.965 ;
        END
        ANTENNAGATEAREA     0.3666 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.730 1.065 1.990 ;
        RECT  0.585 1.700 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.3666 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.645 4.015 1.990 ;
        RECT  3.470 1.645 3.805 1.905 ;
        RECT  3.310 1.645 3.470 2.360 ;
        RECT  2.425 2.200 3.310 2.360 ;
        RECT  2.265 1.645 2.425 2.360 ;
        RECT  2.165 1.645 2.265 1.905 ;
        END
        ANTENNAGATEAREA     0.3666 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.685 1.570 3.095 1.990 ;
        END
        ANTENNAGATEAREA     0.3666 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 -0.250 4.600 0.250 ;
        RECT  1.655 -0.250 1.915 1.060 ;
        RECT  0.895 -0.250 1.655 0.250 ;
        RECT  0.635 -0.250 0.895 1.070 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.785 3.440 4.600 3.940 ;
        RECT  3.525 2.945 3.785 3.940 ;
        RECT  2.085 3.440 3.525 3.940 ;
        RECT  1.825 2.945 2.085 3.940 ;
        RECT  0.385 3.440 1.825 3.940 ;
        RECT  0.125 2.640 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.205 0.605 4.465 0.975 ;
        RECT  3.445 0.605 4.205 0.765 ;
        RECT  3.185 0.605 3.445 0.975 ;
        RECT  2.425 0.605 3.185 0.765 ;
        RECT  2.325 0.605 2.425 1.110 ;
        RECT  2.265 0.605 2.325 1.455 ;
        RECT  2.165 0.850 2.265 1.455 ;
        RECT  1.405 1.295 2.165 1.455 ;
        RECT  1.145 0.850 1.405 1.455 ;
        RECT  0.385 1.295 1.145 1.455 ;
        RECT  0.225 0.850 0.385 1.455 ;
        RECT  0.125 0.850 0.225 1.110 ;
    END
END OAI22X2

MACRO OAI22X1
    CLASS CORE ;
    FOREIGN OAI22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.290 2.635 1.765 ;
        RECT  2.425 1.235 2.585 2.365 ;
        RECT  2.015 1.235 2.425 1.395 ;
        RECT  1.470 2.205 2.425 2.365 ;
        RECT  1.755 0.985 2.015 1.395 ;
        RECT  1.310 2.205 1.470 2.980 ;
        RECT  1.210 2.380 1.310 2.980 ;
        END
        ANTENNADIFFAREA     0.6924 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.405 0.555 1.730 ;
        RECT  0.125 1.405 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.065 1.710 1.165 1.970 ;
        RECT  0.905 1.710 1.065 2.270 ;
        RECT  0.795 2.110 0.905 2.270 ;
        RECT  0.585 2.110 0.795 2.400 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.920 1.580 2.230 2.005 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 1.585 1.735 2.020 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.935 -0.250 2.760 0.250 ;
        RECT  0.675 -0.250 0.935 0.845 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.385 3.440 2.760 3.940 ;
        RECT  2.125 2.545 2.385 3.940 ;
        RECT  0.485 3.440 2.125 3.940 ;
        RECT  0.225 2.580 0.485 3.940 ;
        RECT  0.000 3.440 0.225 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.425 0.795 2.525 1.055 ;
        RECT  2.265 0.645 2.425 1.055 ;
        RECT  1.505 0.645 2.265 0.805 ;
        RECT  1.345 0.645 1.505 1.195 ;
        RECT  1.245 0.935 1.345 1.195 ;
        RECT  0.385 1.035 1.245 1.195 ;
        RECT  0.125 0.935 0.385 1.195 ;
    END
END OAI22X1

MACRO OAI22XL
    CLASS CORE ;
    FOREIGN OAI22XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.755 2.205 2.740 ;
        RECT  2.125 1.290 2.175 2.740 ;
        RECT  2.045 1.125 2.125 2.740 ;
        RECT  2.015 1.125 2.045 1.915 ;
        RECT  1.265 2.580 2.045 2.740 ;
        RECT  1.965 1.125 2.015 1.580 ;
        RECT  1.735 1.125 1.965 1.285 ;
        RECT  1.475 1.025 1.735 1.285 ;
        RECT  1.005 2.580 1.265 2.840 ;
        END
        ANTENNADIFFAREA     0.2888 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.840 0.405 2.400 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.770 0.925 1.930 ;
        RECT  0.635 1.770 0.795 2.400 ;
        RECT  0.585 2.110 0.635 2.400 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.585 2.095 1.865 2.400 ;
        RECT  1.445 2.110 1.585 2.400 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 1.770 1.435 1.930 ;
        RECT  1.105 1.770 1.265 2.400 ;
        RECT  1.045 2.110 1.105 2.400 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 -0.250 2.300 0.250 ;
        RECT  0.625 -0.250 0.785 1.235 ;
        RECT  0.000 -0.250 0.625 0.250 ;
        RECT  0.525 1.075 0.625 1.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 3.440 2.300 3.940 ;
        RECT  1.915 2.945 2.175 3.940 ;
        RECT  0.385 3.440 1.915 3.940 ;
        RECT  0.125 2.725 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.875 0.445 2.135 0.705 ;
        RECT  1.125 0.545 1.875 0.705 ;
        RECT  0.965 0.545 1.125 1.575 ;
        RECT  0.285 1.415 0.965 1.575 ;
        RECT  0.285 0.445 0.385 0.705 ;
        RECT  0.125 0.445 0.285 1.575 ;
    END
END OAI22XL

MACRO OAI211X4
    CLASS CORE ;
    FOREIGN OAI211X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.755 1.010 4.015 2.355 ;
        RECT  3.475 1.010 3.755 1.270 ;
        RECT  3.475 2.095 3.755 2.355 ;
        RECT  3.215 0.635 3.475 1.270 ;
        RECT  3.215 2.095 3.475 3.045 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 1.290 1.405 1.985 ;
        RECT  1.045 1.290 1.145 1.580 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.675 1.605 2.175 2.015 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.405 0.405 1.665 ;
        RECT  0.125 1.405 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 1.760 0.925 2.020 ;
        RECT  0.585 1.470 0.840 2.020 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.985 -0.250 4.140 0.250 ;
        RECT  3.725 -0.250 3.985 0.745 ;
        RECT  2.965 -0.250 3.725 0.250 ;
        RECT  2.705 -0.250 2.965 0.745 ;
        RECT  0.785 -0.250 2.705 0.250 ;
        RECT  0.525 -0.250 0.785 1.195 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.985 3.440 4.140 3.940 ;
        RECT  3.725 2.615 3.985 3.940 ;
        RECT  2.965 3.440 3.725 3.940 ;
        RECT  2.705 2.955 2.965 3.940 ;
        RECT  1.500 3.440 2.705 3.940 ;
        RECT  1.240 3.285 1.500 3.940 ;
        RECT  0.385 3.440 1.240 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.030 1.605 3.305 1.865 ;
        RECT  2.870 0.925 3.030 2.750 ;
        RECT  2.455 0.925 2.870 1.085 ;
        RECT  2.455 2.590 2.870 2.750 ;
        RECT  2.515 1.635 2.615 1.895 ;
        RECT  2.355 1.265 2.515 2.360 ;
        RECT  2.295 0.505 2.455 1.085 ;
        RECT  2.295 2.590 2.455 3.045 ;
        RECT  2.055 1.265 2.355 1.425 ;
        RECT  2.055 2.200 2.355 2.360 ;
        RECT  2.195 0.505 2.295 0.765 ;
        RECT  2.195 2.785 2.295 3.045 ;
        RECT  1.895 1.035 2.055 1.425 ;
        RECT  1.795 2.200 2.055 2.460 ;
        RECT  1.795 1.035 1.895 1.295 ;
        RECT  1.095 2.200 1.795 2.360 ;
        RECT  0.835 2.200 1.095 2.460 ;
    END
END OAI211X4

MACRO OAI211X2
    CLASS CORE ;
    FOREIGN OAI211X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.945 1.925 4.015 2.175 ;
        RECT  3.785 1.420 3.945 2.415 ;
        RECT  3.555 1.420 3.785 1.580 ;
        RECT  3.230 2.255 3.785 2.415 ;
        RECT  3.505 1.290 3.555 1.580 ;
        RECT  3.345 0.810 3.505 1.580 ;
        RECT  2.845 0.810 3.345 0.970 ;
        RECT  2.970 2.255 3.230 3.195 ;
        RECT  2.175 2.255 2.970 2.415 ;
        RECT  2.170 2.255 2.175 2.585 ;
        RECT  1.910 2.255 2.170 2.855 ;
        RECT  0.385 2.580 1.910 2.740 ;
        RECT  0.125 2.265 0.385 2.865 ;
        END
        ANTENNADIFFAREA     1.4640 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.760 3.605 2.020 ;
        RECT  2.635 1.830 3.345 1.990 ;
        RECT  2.455 1.700 2.635 1.990 ;
        RECT  2.195 1.585 2.455 1.990 ;
        END
        ANTENNAGATEAREA     0.3380 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 1.150 3.165 1.650 ;
        END
        ANTENNAGATEAREA     0.3380 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.885 1.375 2.140 ;
        RECT  1.045 1.885 1.255 2.400 ;
        RECT  0.775 1.885 1.045 2.140 ;
        END
        ANTENNAGATEAREA     0.3640 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.815 1.725 1.915 1.985 ;
        RECT  1.655 1.455 1.815 1.985 ;
        RECT  0.555 1.455 1.655 1.615 ;
        RECT  0.335 1.455 0.555 1.715 ;
        RECT  0.295 1.455 0.335 1.990 ;
        RECT  0.125 1.555 0.295 1.990 ;
        END
        ANTENNAGATEAREA     0.3913 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.735 -0.250 4.140 0.250 ;
        RECT  1.475 -0.250 1.735 0.405 ;
        RECT  0.935 -0.250 1.475 0.250 ;
        RECT  0.675 -0.250 0.935 0.405 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.720 3.440 4.140 3.940 ;
        RECT  2.460 2.595 2.720 3.940 ;
        RECT  1.235 3.440 2.460 3.940 ;
        RECT  0.975 2.945 1.235 3.940 ;
        RECT  0.000 3.440 0.975 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.845 0.850 3.945 1.110 ;
        RECT  3.685 0.470 3.845 1.110 ;
        RECT  2.285 0.470 3.685 0.630 ;
        RECT  2.125 0.470 2.285 1.275 ;
        RECT  2.025 0.675 2.125 1.275 ;
        RECT  1.335 1.000 2.025 1.160 ;
        RECT  1.075 0.900 1.335 1.160 ;
        RECT  0.385 1.000 1.075 1.160 ;
        RECT  0.125 0.675 0.385 1.275 ;
    END
END OAI211X2

MACRO OAI211X1
    CLASS CORE ;
    FOREIGN OAI211X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.170 0.695 2.175 2.360 ;
        RECT  1.910 0.685 2.170 2.620 ;
        RECT  1.255 2.360 1.910 2.570 ;
        RECT  1.045 2.360 1.255 2.810 ;
        RECT  0.955 2.360 1.045 2.620 ;
        END
        ANTENNADIFFAREA     0.7376 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.700 1.715 2.090 ;
        END
        ANTENNAGATEAREA     0.1690 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 2.850 2.175 3.220 ;
        RECT  1.825 2.850 1.965 3.205 ;
        END
        ANTENNAGATEAREA     0.1690 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.520 0.360 2.070 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.430 1.035 1.815 ;
        RECT  0.585 1.290 0.835 1.815 ;
        END
        ANTENNAGATEAREA     0.1820 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.935 -0.250 2.300 0.250 ;
        RECT  0.675 -0.250 0.935 0.405 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.615 3.440 2.300 3.940 ;
        RECT  1.355 3.285 1.615 3.940 ;
        RECT  0.385 3.440 1.355 3.940 ;
        RECT  0.125 2.420 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.075 0.860 1.335 1.120 ;
        RECT  0.385 0.860 1.075 1.020 ;
        RECT  0.125 0.675 0.385 1.275 ;
    END
END OAI211X1

MACRO OAI211XL
    CLASS CORE ;
    FOREIGN OAI211XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.165 1.105 2.175 2.620 ;
        RECT  1.965 0.935 2.165 2.620 ;
        RECT  1.905 0.935 1.965 1.195 ;
        RECT  1.915 2.325 1.965 2.620 ;
        RECT  1.255 2.325 1.915 2.520 ;
        RECT  1.045 2.325 1.255 2.810 ;
        RECT  1.035 2.325 1.045 2.725 ;
        RECT  0.945 2.465 1.035 2.725 ;
        END
        ANTENNADIFFAREA     0.4182 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.700 1.715 1.990 ;
        RECT  1.260 1.715 1.505 1.975 ;
        END
        ANTENNAGATEAREA     0.0910 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 2.830 2.175 3.220 ;
        RECT  1.725 2.830 1.965 3.055 ;
        END
        ANTENNAGATEAREA     0.0910 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.525 0.360 2.130 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.635 1.035 1.895 ;
        RECT  0.830 1.355 0.835 1.895 ;
        RECT  0.645 1.290 0.830 1.895 ;
        RECT  0.585 1.290 0.645 1.765 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 -0.250 2.300 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 3.440 2.300 3.940 ;
        RECT  1.375 3.285 1.635 3.940 ;
        RECT  0.385 3.440 1.375 3.940 ;
        RECT  0.125 2.625 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.085 0.910 1.345 1.170 ;
        RECT  0.385 0.910 1.085 1.070 ;
        RECT  0.125 0.910 0.385 1.170 ;
    END
END OAI211XL

MACRO OAI21X4
    CLASS CORE ;
    FOREIGN OAI21X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 0.640 4.935 2.335 ;
        RECT  4.725 0.640 4.885 2.390 ;
        RECT  4.675 0.640 4.725 1.520 ;
        RECT  4.065 2.230 4.725 2.390 ;
        RECT  3.915 1.360 4.675 1.520 ;
        RECT  3.905 2.230 4.065 2.735 ;
        RECT  3.755 1.035 3.915 1.520 ;
        RECT  3.805 2.455 3.905 2.735 ;
        RECT  3.045 2.455 3.805 2.615 ;
        RECT  3.655 1.035 3.755 1.295 ;
        RECT  2.610 2.455 3.045 3.055 ;
        RECT  1.305 2.455 2.610 2.615 ;
        RECT  1.045 2.455 1.305 3.055 ;
        END
        ANTENNADIFFAREA     1.7037 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.740 4.090 2.000 ;
        RECT  3.805 1.700 4.015 2.000 ;
        RECT  3.490 1.740 3.805 2.000 ;
        END
        ANTENNAGATEAREA     0.6318 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.025 1.615 2.285 1.875 ;
        RECT  1.475 1.615 2.025 1.775 ;
        RECT  1.315 1.475 1.475 1.775 ;
        RECT  0.655 1.475 1.315 1.635 ;
        RECT  0.395 1.475 0.655 1.770 ;
        RECT  0.335 1.610 0.395 1.770 ;
        RECT  0.125 1.610 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.7371 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 1.715 3.075 1.975 ;
        RECT  2.815 1.715 2.975 2.270 ;
        RECT  1.135 2.110 2.815 2.270 ;
        RECT  0.875 1.815 1.135 2.270 ;
        RECT  0.795 2.110 0.875 2.270 ;
        RECT  0.585 2.110 0.795 2.400 ;
        END
        ANTENNAGATEAREA     0.7306 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.005 -0.250 5.060 0.250 ;
        RECT  2.745 -0.250 3.005 0.405 ;
        RECT  1.915 -0.250 2.745 0.250 ;
        RECT  1.655 -0.250 1.915 0.955 ;
        RECT  0.895 -0.250 1.655 0.250 ;
        RECT  0.635 -0.250 0.895 0.840 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 3.440 5.060 3.940 ;
        RECT  4.315 2.725 4.575 3.940 ;
        RECT  3.555 3.440 4.315 3.940 ;
        RECT  3.295 2.950 3.555 3.940 ;
        RECT  2.185 3.440 3.295 3.940 ;
        RECT  1.925 2.955 2.185 3.940 ;
        RECT  0.485 3.440 1.925 3.940 ;
        RECT  0.225 2.615 0.485 3.940 ;
        RECT  0.000 3.440 0.225 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.165 0.565 4.425 1.165 ;
        RECT  3.405 0.695 4.165 0.855 ;
        RECT  3.145 0.695 3.405 1.070 ;
        RECT  2.425 0.910 3.145 1.070 ;
        RECT  2.165 0.810 2.425 1.410 ;
        RECT  1.405 1.135 2.165 1.295 ;
        RECT  1.145 0.640 1.405 1.295 ;
        RECT  0.385 1.135 1.145 1.295 ;
        RECT  0.125 0.640 0.385 1.295 ;
    END
END OAI21X4

MACRO OAI21X2
    CLASS CORE ;
    FOREIGN OAI21X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.015 1.290 3.095 1.765 ;
        RECT  2.910 0.945 3.015 2.330 ;
        RECT  2.855 0.945 2.910 2.335 ;
        RECT  2.755 0.945 2.855 1.205 ;
        RECT  2.765 2.170 2.855 2.335 ;
        RECT  2.505 2.170 2.765 2.770 ;
        RECT  2.425 2.230 2.505 2.585 ;
        RECT  1.305 2.230 2.425 2.390 ;
        RECT  1.045 2.230 1.305 2.830 ;
        END
        ANTENNADIFFAREA     0.7828 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.340 1.510 2.675 1.990 ;
        END
        ANTENNAGATEAREA     0.3172 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.855 1.665 1.955 1.925 ;
        RECT  1.695 1.450 1.855 1.925 ;
        RECT  0.455 1.450 1.695 1.610 ;
        RECT  0.385 1.450 0.455 1.770 ;
        RECT  0.125 1.450 0.385 1.990 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.975 1.790 1.235 2.050 ;
        RECT  0.795 1.890 0.975 2.050 ;
        RECT  0.635 1.890 0.795 2.400 ;
        RECT  0.585 2.110 0.635 2.400 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 -0.250 3.680 0.250 ;
        RECT  1.695 -0.250 1.955 0.795 ;
        RECT  0.895 -0.250 1.695 0.250 ;
        RECT  0.635 -0.250 0.895 0.930 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.305 3.440 3.680 3.940 ;
        RECT  3.045 2.555 3.305 3.940 ;
        RECT  2.225 3.440 3.045 3.940 ;
        RECT  1.965 2.895 2.225 3.940 ;
        RECT  0.385 3.440 1.965 3.940 ;
        RECT  0.125 2.555 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.265 0.605 3.525 0.930 ;
        RECT  2.505 0.605 3.265 0.765 ;
        RECT  2.405 0.605 2.505 0.930 ;
        RECT  2.245 0.605 2.405 1.270 ;
        RECT  1.405 1.110 2.245 1.270 ;
        RECT  1.145 0.950 1.405 1.270 ;
        RECT  0.385 1.110 1.145 1.270 ;
        RECT  0.125 0.950 0.385 1.270 ;
    END
END OAI21X2

MACRO OAI21X1
    CLASS CORE ;
    FOREIGN OAI21X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.990 1.010 2.175 2.400 ;
        RECT  1.965 0.910 1.990 2.400 ;
        RECT  1.655 0.910 1.965 1.170 ;
        RECT  1.275 2.230 1.965 2.390 ;
        RECT  1.015 2.230 1.275 2.830 ;
        END
        ANTENNADIFFAREA     0.4864 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.355 1.635 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.1586 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.145 1.510 0.405 1.990 ;
        RECT  0.125 1.700 0.145 1.990 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.510 1.035 1.770 ;
        RECT  0.635 1.510 0.795 2.400 ;
        RECT  0.585 1.925 0.635 2.400 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 -0.250 2.300 0.250 ;
        RECT  0.635 -0.250 0.895 0.990 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 3.440 2.300 3.940 ;
        RECT  1.525 2.570 1.785 3.940 ;
        RECT  0.385 3.440 1.525 3.940 ;
        RECT  0.125 2.330 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.145 0.910 1.405 1.330 ;
        RECT  0.385 1.170 1.145 1.330 ;
        RECT  0.125 0.925 0.385 1.330 ;
    END
END OAI21X1

MACRO OAI21XL
    CLASS CORE ;
    FOREIGN OAI21XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.695 0.695 1.715 1.990 ;
        RECT  1.665 0.445 1.695 1.990 ;
        RECT  1.505 0.445 1.665 2.240 ;
        RECT  1.435 0.445 1.505 0.705 ;
        RECT  1.235 2.080 1.505 2.240 ;
        RECT  0.975 2.080 1.235 2.340 ;
        END
        ANTENNADIFFAREA     0.3680 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 2.520 1.405 2.865 ;
        RECT  0.975 2.520 1.145 2.860 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.550 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.470 1.035 1.730 ;
        RECT  0.775 1.470 0.795 2.400 ;
        RECT  0.635 1.570 0.775 2.400 ;
        RECT  0.585 1.925 0.635 2.400 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 -0.250 1.840 0.250 ;
        RECT  0.635 -0.250 0.895 0.405 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 3.440 1.840 3.940 ;
        RECT  1.375 3.285 1.635 3.940 ;
        RECT  0.385 3.440 1.375 3.940 ;
        RECT  0.125 2.230 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.035 1.030 1.295 1.290 ;
        RECT  0.385 1.030 1.035 1.190 ;
        RECT  0.225 0.445 0.385 1.190 ;
        RECT  0.125 0.445 0.225 0.705 ;
    END
END OAI21XL

MACRO OR4X8
    CLASS CORE ;
    FOREIGN OR4X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.180 1.105 7.235 2.585 ;
        RECT  6.920 0.635 7.180 2.965 ;
        RECT  6.160 0.975 6.920 2.115 ;
        RECT  6.105 0.635 6.160 2.965 ;
        RECT  5.900 0.635 6.105 1.235 ;
        RECT  5.900 1.855 6.105 2.965 ;
        END
        ANTENNADIFFAREA     1.5812 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.275 1.745 5.375 2.005 ;
        RECT  5.115 1.745 5.275 2.685 ;
        RECT  2.175 2.525 5.115 2.685 ;
        RECT  2.015 1.805 2.175 2.685 ;
        RECT  1.965 1.805 2.015 2.400 ;
        RECT  1.700 1.805 1.965 1.965 ;
        END
        ANTENNAGATEAREA     0.5863 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.685 1.405 4.845 2.345 ;
        RECT  2.635 2.185 4.685 2.345 ;
        RECT  2.475 1.465 2.635 2.345 ;
        RECT  2.425 1.465 2.475 1.990 ;
        RECT  1.180 1.465 2.425 1.625 ;
        END
        ANTENNAGATEAREA     0.5863 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.315 1.290 4.475 1.765 ;
        RECT  4.155 1.290 4.315 2.005 ;
        RECT  3.095 1.845 4.155 2.005 ;
        RECT  3.020 1.515 3.095 2.005 ;
        RECT  2.860 1.125 3.020 2.005 ;
        RECT  1.130 1.125 2.860 1.285 ;
        RECT  0.870 0.935 1.130 1.285 ;
        END
        ANTENNAGATEAREA     0.5863 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.290 3.820 1.665 ;
        END
        ANTENNAGATEAREA     0.5863 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.690 -0.250 7.820 0.250 ;
        RECT  7.430 -0.250 7.690 1.090 ;
        RECT  6.670 -0.250 7.430 0.250 ;
        RECT  6.410 -0.250 6.670 0.755 ;
        RECT  5.650 -0.250 6.410 0.250 ;
        RECT  5.390 -0.250 5.650 0.750 ;
        RECT  4.560 -0.250 5.390 0.250 ;
        RECT  4.300 -0.250 4.560 0.405 ;
        RECT  3.760 -0.250 4.300 0.250 ;
        RECT  3.500 -0.250 3.760 0.405 ;
        RECT  2.670 -0.250 3.500 0.250 ;
        RECT  2.410 -0.250 2.670 0.605 ;
        RECT  1.620 -0.250 2.410 0.250 ;
        RECT  1.360 -0.250 1.620 0.945 ;
        RECT  0.000 -0.250 1.360 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.690 3.440 7.820 3.940 ;
        RECT  7.430 2.075 7.690 3.940 ;
        RECT  6.670 3.440 7.430 3.940 ;
        RECT  6.410 2.415 6.670 3.940 ;
        RECT  5.470 3.440 6.410 3.940 ;
        RECT  5.210 3.285 5.470 3.940 ;
        RECT  2.000 3.440 5.210 3.940 ;
        RECT  1.740 3.285 2.000 3.940 ;
        RECT  0.000 3.440 1.740 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.720 1.415 5.875 1.675 ;
        RECT  5.560 0.930 5.720 3.025 ;
        RECT  5.110 0.930 5.560 1.090 ;
        RECT  3.905 2.865 5.560 3.025 ;
        RECT  4.850 0.830 5.110 1.090 ;
        RECT  4.160 0.930 4.850 1.090 ;
        RECT  3.900 0.785 4.160 1.090 ;
        RECT  3.305 2.865 3.905 3.125 ;
        RECT  3.210 0.785 3.900 0.945 ;
        RECT  0.480 2.865 3.305 3.025 ;
        RECT  2.950 0.685 3.210 0.945 ;
        RECT  2.130 0.785 2.950 0.945 ;
        RECT  1.870 0.685 2.130 0.945 ;
        RECT  0.220 2.125 0.480 3.065 ;
    END
END OR4X8

MACRO OR4X6
    CLASS CORE ;
    FOREIGN OR4X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.590 0.635 5.855 1.290 ;
        RECT  5.850 1.855 5.855 2.585 ;
        RECT  5.590 1.855 5.850 2.965 ;
        RECT  5.395 0.975 5.590 1.290 ;
        RECT  5.395 1.855 5.590 2.155 ;
        RECT  4.830 0.975 5.395 2.155 ;
        RECT  4.725 0.635 4.830 2.965 ;
        RECT  4.570 0.635 4.725 1.235 ;
        RECT  4.570 1.855 4.725 2.965 ;
        END
        ANTENNADIFFAREA     1.4584 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.675 4.045 1.935 ;
        RECT  3.945 1.675 4.015 2.175 ;
        RECT  3.785 1.675 3.945 2.605 ;
        RECT  0.915 2.445 3.785 2.605 ;
        RECT  0.795 1.865 0.915 2.605 ;
        RECT  0.755 1.290 0.795 2.605 ;
        RECT  0.635 1.290 0.755 2.025 ;
        RECT  0.585 1.290 0.635 1.765 ;
        RECT  0.490 1.315 0.585 1.575 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.315 3.565 1.575 ;
        RECT  3.465 1.315 3.555 1.765 ;
        RECT  3.305 1.315 3.465 2.260 ;
        RECT  1.255 2.100 3.305 2.260 ;
        RECT  1.095 1.290 1.255 2.260 ;
        RECT  0.980 1.290 1.095 1.580 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.985 1.290 3.095 1.580 ;
        RECT  2.885 1.290 2.985 1.920 ;
        RECT  2.825 1.315 2.885 1.920 ;
        RECT  1.715 1.760 2.825 1.920 ;
        RECT  1.555 1.360 1.715 1.920 ;
        RECT  1.455 1.360 1.555 1.620 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 1.290 2.635 1.580 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.340 -0.250 5.980 0.250 ;
        RECT  5.080 -0.250 5.340 0.755 ;
        RECT  4.320 -0.250 5.080 0.250 ;
        RECT  4.060 -0.250 4.320 0.750 ;
        RECT  3.230 -0.250 4.060 0.250 ;
        RECT  2.970 -0.250 3.230 0.405 ;
        RECT  2.430 -0.250 2.970 0.250 ;
        RECT  2.170 -0.250 2.430 0.405 ;
        RECT  1.480 -0.250 2.170 0.250 ;
        RECT  1.220 -0.250 1.480 0.405 ;
        RECT  0.420 -0.250 1.220 0.250 ;
        RECT  0.160 -0.250 0.420 1.035 ;
        RECT  0.000 -0.250 0.160 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.340 3.440 5.980 3.940 ;
        RECT  5.080 2.415 5.340 3.940 ;
        RECT  4.140 3.440 5.080 3.940 ;
        RECT  3.880 3.285 4.140 3.940 ;
        RECT  0.570 3.440 3.880 3.940 ;
        RECT  0.310 2.275 0.570 3.940 ;
        RECT  0.000 3.440 0.310 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.390 1.415 4.545 1.675 ;
        RECT  4.230 0.930 4.390 2.945 ;
        RECT  3.780 0.930 4.230 1.090 ;
        RECT  2.535 2.785 4.230 2.945 ;
        RECT  3.520 0.830 3.780 1.090 ;
        RECT  2.830 0.930 3.520 1.090 ;
        RECT  2.570 0.830 2.830 1.090 ;
        RECT  2.565 0.880 2.570 1.090 ;
        RECT  1.880 0.930 2.565 1.090 ;
        RECT  1.935 2.785 2.535 3.045 ;
        RECT  1.620 0.830 1.880 1.090 ;
        RECT  0.930 0.930 1.620 1.090 ;
        RECT  0.670 0.830 0.930 1.090 ;
    END
END OR4X6

MACRO OR4X4
    CLASS CORE ;
    FOREIGN OR4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.215 0.940 4.475 2.365 ;
        RECT  3.945 0.940 4.215 1.200 ;
        RECT  4.015 2.105 4.215 2.365 ;
        RECT  3.945 2.105 4.015 2.585 ;
        RECT  3.685 0.600 3.945 1.200 ;
        RECT  3.685 2.105 3.945 3.095 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.995 1.925 3.095 2.185 ;
        RECT  2.835 1.925 2.995 2.630 ;
        RECT  0.385 2.470 2.835 2.630 ;
        RECT  0.225 1.740 0.385 2.630 ;
        RECT  0.125 1.740 0.225 2.405 ;
        END
        ANTENNAGATEAREA     0.3289 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 1.445 2.785 1.705 ;
        RECT  2.525 1.445 2.610 1.765 ;
        RECT  2.515 1.545 2.525 1.765 ;
        RECT  2.355 1.545 2.515 2.290 ;
        RECT  0.795 2.130 2.355 2.290 ;
        RECT  0.635 1.360 0.795 2.290 ;
        RECT  0.585 1.360 0.635 1.990 ;
        RECT  0.545 1.360 0.585 1.520 ;
        RECT  0.285 1.260 0.545 1.520 ;
        END
        ANTENNAGATEAREA     0.3289 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.165 1.290 2.175 1.580 ;
        RECT  2.065 1.280 2.165 1.580 ;
        RECT  1.905 1.280 2.065 1.950 ;
        RECT  1.135 1.790 1.905 1.950 ;
        RECT  0.975 1.000 1.135 1.950 ;
        RECT  0.765 1.000 0.975 1.160 ;
        END
        ANTENNAGATEAREA     0.3289 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.560 1.280 1.715 1.610 ;
        RECT  1.315 1.020 1.560 1.610 ;
        END
        ANTENNAGATEAREA     0.3289 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.455 -0.250 4.600 0.250 ;
        RECT  4.195 -0.250 4.455 0.755 ;
        RECT  3.435 -0.250 4.195 0.250 ;
        RECT  3.175 -0.250 3.435 0.755 ;
        RECT  2.415 -0.250 3.175 0.250 ;
        RECT  2.155 -0.250 2.415 0.755 ;
        RECT  1.395 -0.250 2.155 0.250 ;
        RECT  1.135 -0.250 1.395 0.755 ;
        RECT  0.000 -0.250 1.135 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.455 3.440 4.600 3.940 ;
        RECT  4.195 2.545 4.455 3.940 ;
        RECT  3.320 3.440 4.195 3.940 ;
        RECT  3.060 3.285 3.320 3.940 ;
        RECT  0.385 3.440 3.060 3.940 ;
        RECT  0.125 2.810 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.435 1.555 3.775 1.815 ;
        RECT  3.275 0.935 3.435 2.970 ;
        RECT  2.925 0.935 3.275 1.095 ;
        RECT  1.565 2.810 3.275 2.970 ;
        RECT  2.665 0.495 2.925 1.095 ;
        RECT  1.905 0.935 2.665 1.095 ;
        RECT  1.745 0.545 1.905 1.095 ;
        RECT  1.645 0.545 1.745 0.805 ;
    END
END OR4X4

MACRO OR4X2
    CLASS CORE ;
    FOREIGN OR4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 0.490 3.095 3.055 ;
        RECT  2.835 0.490 2.935 1.090 ;
        RECT  2.885 2.110 2.935 3.055 ;
        RECT  2.835 2.115 2.885 3.055 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 2.110 2.635 2.400 ;
        RECT  2.425 1.860 2.585 2.400 ;
        RECT  2.315 1.860 2.425 2.020 ;
        RECT  2.055 1.760 2.315 2.020 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.875 1.280 2.005 1.580 ;
        RECT  1.715 1.280 1.875 1.925 ;
        RECT  1.505 1.700 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.260 1.535 1.520 ;
        RECT  0.975 1.260 1.255 1.580 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.915 1.760 1.175 2.020 ;
        RECT  0.795 1.760 0.915 1.990 ;
        RECT  0.770 1.290 0.795 1.990 ;
        RECT  0.585 1.290 0.770 1.920 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 -0.250 3.220 0.250 ;
        RECT  2.285 -0.250 2.545 0.405 ;
        RECT  1.745 -0.250 2.285 0.250 ;
        RECT  1.485 -0.250 1.745 0.405 ;
        RECT  0.655 -0.250 1.485 0.250 ;
        RECT  0.395 -0.250 0.655 0.405 ;
        RECT  0.000 -0.250 0.395 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 3.440 3.220 3.940 ;
        RECT  2.325 2.595 2.585 3.940 ;
        RECT  0.000 3.440 2.325 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.655 1.400 2.755 1.660 ;
        RECT  2.495 0.920 2.655 1.660 ;
        RECT  2.145 0.920 2.495 1.080 ;
        RECT  1.885 0.820 2.145 1.080 ;
        RECT  1.195 0.920 1.885 1.080 ;
        RECT  0.935 0.820 1.195 1.080 ;
        RECT  0.745 2.275 1.005 2.875 ;
        RECT  0.405 0.920 0.935 1.080 ;
        RECT  0.405 2.275 0.745 2.435 ;
        RECT  0.245 0.920 0.405 2.435 ;
    END
END OR4X2

MACRO OR4X1
    CLASS CORE ;
    FOREIGN OR4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 0.895 2.635 3.020 ;
        RECT  2.425 0.895 2.475 1.580 ;
        RECT  2.375 2.420 2.475 3.020 ;
        RECT  2.375 0.895 2.425 1.155 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 0.880 2.175 1.170 ;
        RECT  1.965 0.880 1.985 1.610 ;
        RECT  1.825 0.945 1.965 1.610 ;
        RECT  1.775 1.350 1.825 1.610 ;
        END
        ANTENNAGATEAREA     0.0806 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.095 1.350 1.255 2.400 ;
        RECT  1.045 1.925 1.095 2.400 ;
        END
        ANTENNAGATEAREA     0.0806 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.455 1.290 0.795 1.920 ;
        END
        ANTENNAGATEAREA     0.0806 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.140 0.765 2.400 ;
        RECT  0.125 2.110 0.335 2.400 ;
        END
        ANTENNAGATEAREA     0.0806 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 -0.250 2.760 0.250 ;
        RECT  1.975 -0.250 2.235 0.405 ;
        RECT  1.205 -0.250 1.975 0.250 ;
        RECT  0.945 -0.250 1.205 0.405 ;
        RECT  0.545 -0.250 0.945 0.250 ;
        RECT  0.285 -0.250 0.545 0.405 ;
        RECT  0.000 -0.250 0.285 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 3.440 2.760 3.940 ;
        RECT  1.865 2.420 2.125 3.940 ;
        RECT  0.000 3.440 1.865 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.595 1.865 2.295 2.125 ;
        RECT  1.595 0.910 1.645 1.170 ;
        RECT  1.435 0.910 1.595 2.790 ;
        RECT  1.385 0.910 1.435 1.170 ;
        RECT  0.595 2.630 1.435 2.790 ;
        RECT  0.615 0.950 1.385 1.110 ;
        RECT  0.355 0.815 0.615 1.110 ;
        RECT  0.335 2.630 0.595 2.890 ;
    END
END OR4X1

MACRO OR4XL
    CLASS CORE ;
    FOREIGN OR4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.630 0.695 2.635 2.640 ;
        RECT  2.600 0.695 2.630 2.900 ;
        RECT  2.370 0.550 2.600 2.900 ;
        RECT  2.340 0.550 2.370 0.810 ;
        END
        ANTENNADIFFAREA     0.3296 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.085 1.290 2.175 1.765 ;
        RECT  1.925 1.290 2.085 2.000 ;
        RECT  1.825 1.740 1.925 2.000 ;
        END
        ANTENNAGATEAREA     0.0767 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.340 1.305 1.600 ;
        RECT  1.045 1.340 1.255 2.400 ;
        END
        ANTENNAGATEAREA     0.0767 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.300 0.815 1.910 ;
        RECT  0.585 1.290 0.795 1.910 ;
        RECT  0.555 1.300 0.585 1.910 ;
        END
        ANTENNAGATEAREA     0.0767 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 2.110 0.590 2.455 ;
        END
        ANTENNAGATEAREA     0.0767 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.085 -0.250 2.760 0.250 ;
        RECT  1.825 -0.250 2.085 0.405 ;
        RECT  1.055 -0.250 1.825 0.250 ;
        RECT  0.355 -0.250 1.055 0.405 ;
        RECT  0.000 -0.250 0.355 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.090 3.440 2.760 3.940 ;
        RECT  1.830 2.665 2.090 3.940 ;
        RECT  0.000 3.440 1.830 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.645 2.225 2.175 2.485 ;
        RECT  1.485 0.900 1.645 2.900 ;
        RECT  1.385 0.900 1.485 1.160 ;
        RECT  0.595 2.740 1.485 2.900 ;
        RECT  0.615 0.945 1.385 1.105 ;
        RECT  0.355 0.815 0.615 1.105 ;
        RECT  0.335 2.740 0.595 3.000 ;
    END
END OR4XL

MACRO OR3X8
    CLASS CORE ;
    FOREIGN OR3X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 0.925 5.870 1.405 ;
        RECT  5.805 0.580 5.855 2.585 ;
        RECT  5.545 0.580 5.805 3.065 ;
        RECT  5.185 0.925 5.545 2.595 ;
        RECT  4.850 0.925 5.185 1.405 ;
        RECT  4.785 2.005 5.185 2.595 ;
        RECT  4.575 0.580 4.850 1.405 ;
        RECT  4.640 2.005 4.785 3.135 ;
        RECT  4.525 2.435 4.640 3.135 ;
        END
        ANTENNADIFFAREA     1.6112 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.895 1.035 4.055 1.780 ;
        RECT  3.805 1.035 3.895 1.355 ;
        RECT  1.860 1.035 3.805 1.195 ;
        RECT  1.700 1.035 1.860 1.580 ;
        RECT  1.505 1.290 1.700 1.580 ;
        END
        ANTENNAGATEAREA     0.5577 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.520 1.620 3.620 1.880 ;
        RECT  3.360 1.380 3.520 1.880 ;
        RECT  2.540 1.380 3.360 1.540 ;
        RECT  2.440 1.380 2.540 1.570 ;
        RECT  2.280 1.380 2.440 1.940 ;
        RECT  1.255 1.780 2.280 1.940 ;
        RECT  1.045 1.290 1.255 1.940 ;
        RECT  0.780 1.680 1.045 1.940 ;
        END
        ANTENNAGATEAREA     0.5577 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.985 1.720 3.105 1.880 ;
        RECT  2.825 1.720 2.985 2.280 ;
        RECT  0.515 2.120 2.825 2.280 ;
        RECT  0.355 1.635 0.515 2.280 ;
        RECT  0.255 1.635 0.355 1.990 ;
        RECT  0.125 1.700 0.255 1.990 ;
        END
        ANTENNAGATEAREA     0.5577 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 -0.250 6.440 0.250 ;
        RECT  6.055 -0.250 6.315 1.180 ;
        RECT  5.295 -0.250 6.055 0.250 ;
        RECT  5.035 -0.250 5.295 0.705 ;
        RECT  4.190 -0.250 5.035 0.250 ;
        RECT  3.930 -0.250 4.190 0.405 ;
        RECT  3.090 -0.250 3.930 0.250 ;
        RECT  2.830 -0.250 3.090 0.405 ;
        RECT  1.990 -0.250 2.830 0.250 ;
        RECT  1.730 -0.250 1.990 0.405 ;
        RECT  0.930 -0.250 1.730 0.250 ;
        RECT  0.670 -0.250 0.930 1.000 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 3.440 6.440 3.940 ;
        RECT  6.055 2.220 6.315 3.940 ;
        RECT  5.295 3.440 6.055 3.940 ;
        RECT  5.035 2.855 5.295 3.940 ;
        RECT  4.275 3.440 5.035 3.940 ;
        RECT  4.015 2.420 4.275 3.940 ;
        RECT  1.695 3.440 4.015 3.940 ;
        RECT  1.435 2.810 1.695 3.940 ;
        RECT  0.000 3.440 1.435 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.395 1.620 4.955 1.780 ;
        RECT  4.235 0.695 4.395 2.230 ;
        RECT  3.640 0.695 4.235 0.855 ;
        RECT  3.790 2.070 4.235 2.230 ;
        RECT  3.630 2.070 3.790 2.620 ;
        RECT  3.380 0.595 3.640 0.855 ;
        RECT  2.965 2.460 3.630 2.620 ;
        RECT  2.540 0.695 3.380 0.855 ;
        RECT  2.705 2.460 2.965 2.720 ;
        RECT  0.385 2.460 2.705 2.620 ;
        RECT  2.280 0.595 2.540 0.855 ;
        RECT  1.440 0.695 2.280 0.855 ;
        RECT  1.180 0.670 1.440 0.930 ;
        RECT  0.125 2.460 0.385 2.720 ;
    END
END OR3X8

MACRO OR3X6
    CLASS CORE ;
    FOREIGN OR3X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.460 0.695 4.475 2.995 ;
        RECT  4.210 0.695 4.460 3.020 ;
        RECT  4.200 0.965 4.210 3.020 ;
        RECT  3.450 0.965 4.200 2.400 ;
        RECT  3.390 0.695 3.450 2.400 ;
        RECT  3.330 0.695 3.390 2.985 ;
        RECT  3.190 0.695 3.330 1.325 ;
        RECT  3.230 2.040 3.330 2.985 ;
        END
        ANTENNADIFFAREA     1.4333 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 1.525 2.635 2.365 ;
        RECT  0.610 2.205 2.475 2.365 ;
        RECT  0.455 2.175 0.610 2.365 ;
        RECT  0.455 1.515 0.555 1.775 ;
        RECT  0.295 1.515 0.455 2.365 ;
        RECT  0.125 1.700 0.295 1.990 ;
        END
        ANTENNAGATEAREA     0.4056 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 1.425 2.135 2.020 ;
        RECT  1.040 1.860 1.975 2.020 ;
        RECT  0.895 1.300 1.040 2.020 ;
        RECT  0.880 0.880 0.895 2.020 ;
        RECT  0.735 0.880 0.880 1.560 ;
        RECT  0.585 0.880 0.735 1.170 ;
        END
        ANTENNAGATEAREA     0.4056 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.305 1.290 1.765 1.635 ;
        END
        ANTENNAGATEAREA     0.4056 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.960 -0.250 4.600 0.250 ;
        RECT  3.700 -0.250 3.960 0.755 ;
        RECT  2.905 -0.250 3.700 0.250 ;
        RECT  2.645 -0.250 2.905 0.805 ;
        RECT  1.845 -0.250 2.645 0.250 ;
        RECT  1.585 -0.250 1.845 0.755 ;
        RECT  0.000 -0.250 1.585 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.950 3.440 4.600 3.940 ;
        RECT  3.690 2.610 3.950 3.940 ;
        RECT  2.930 3.440 3.690 3.940 ;
        RECT  2.670 2.930 2.930 3.940 ;
        RECT  0.385 3.440 2.670 3.940 ;
        RECT  0.125 2.555 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.980 1.530 3.120 1.810 ;
        RECT  2.820 1.010 2.980 2.715 ;
        RECT  2.355 1.010 2.820 1.170 ;
        RECT  1.655 2.555 2.820 2.715 ;
        RECT  2.095 0.570 2.355 1.170 ;
        RECT  1.335 0.950 2.095 1.110 ;
        RECT  1.395 2.555 1.655 3.155 ;
        RECT  1.075 0.510 1.335 1.110 ;
    END
END OR3X6

MACRO OR3X4
    CLASS CORE ;
    FOREIGN OR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 1.290 3.555 1.990 ;
        RECT  3.455 1.045 3.460 1.990 ;
        RECT  3.215 1.045 3.455 2.300 ;
        RECT  3.095 1.045 3.215 1.285 ;
        RECT  3.095 2.060 3.215 2.300 ;
        RECT  3.090 0.695 3.095 1.285 ;
        RECT  2.835 2.060 3.095 3.000 ;
        RECT  2.835 0.615 3.090 1.285 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.155 1.525 2.315 2.050 ;
        RECT  1.740 1.890 2.155 2.050 ;
        RECT  1.580 1.890 1.740 2.400 ;
        RECT  0.610 2.240 1.580 2.400 ;
        RECT  0.445 2.110 0.610 2.400 ;
        RECT  0.185 1.790 0.445 2.400 ;
        RECT  0.125 1.925 0.185 2.400 ;
        END
        ANTENNAGATEAREA     0.3029 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.595 1.350 1.855 1.610 ;
        RECT  0.795 1.350 1.595 1.510 ;
        RECT  0.670 1.290 0.795 1.580 ;
        RECT  0.585 1.255 0.670 1.580 ;
        RECT  0.510 1.255 0.585 1.515 ;
        END
        ANTENNAGATEAREA     0.3029 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.985 1.700 1.395 2.010 ;
        END
        ANTENNAGATEAREA     0.3029 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 -0.250 3.680 0.250 ;
        RECT  3.295 -0.250 3.555 0.805 ;
        RECT  2.535 -0.250 3.295 0.250 ;
        RECT  2.275 -0.250 2.535 0.805 ;
        RECT  1.515 -0.250 2.275 0.250 ;
        RECT  1.255 -0.250 1.515 0.755 ;
        RECT  0.000 -0.250 1.255 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 3.440 3.680 3.940 ;
        RECT  3.295 2.555 3.555 3.940 ;
        RECT  2.535 3.440 3.295 3.940 ;
        RECT  2.275 2.585 2.535 3.940 ;
        RECT  0.385 3.440 2.275 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.655 1.545 2.935 1.805 ;
        RECT  2.495 0.995 2.655 2.400 ;
        RECT  2.025 0.995 2.495 1.155 ;
        RECT  2.095 2.240 2.495 2.400 ;
        RECT  1.935 2.240 2.095 2.815 ;
        RECT  1.765 0.555 2.025 1.155 ;
        RECT  1.405 2.655 1.935 2.815 ;
        RECT  1.010 0.940 1.765 1.100 ;
        RECT  1.145 2.655 1.405 2.915 ;
        RECT  0.850 0.695 1.010 1.100 ;
        RECT  0.745 0.695 0.850 0.955 ;
    END
END OR3X4

MACRO OR3X2
    CLASS CORE ;
    FOREIGN OR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.105 2.635 2.585 ;
        RECT  2.455 0.640 2.585 2.585 ;
        RECT  2.385 0.640 2.455 3.080 ;
        RECT  2.325 0.640 2.385 1.240 ;
        RECT  2.175 2.140 2.385 3.080 ;
        END
        ANTENNADIFFAREA     0.7720 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.605 2.080 1.715 2.415 ;
        RECT  1.345 1.840 1.605 2.415 ;
        END
        ANTENNAGATEAREA     0.1495 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.330 1.580 1.610 ;
        RECT  1.045 1.290 1.255 1.610 ;
        RECT  1.010 1.350 1.045 1.610 ;
        END
        ANTENNAGATEAREA     0.1495 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.635 0.415 2.065 ;
        END
        ANTENNAGATEAREA     0.1495 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 -0.250 2.760 0.250 ;
        RECT  1.775 -0.250 2.035 0.745 ;
        RECT  0.935 -0.250 1.775 0.250 ;
        RECT  0.675 -0.250 0.935 0.745 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.845 3.440 2.760 3.940 ;
        RECT  1.585 2.710 1.845 3.940 ;
        RECT  0.000 3.440 1.585 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.050 1.575 2.150 1.835 ;
        RECT  1.890 0.925 2.050 1.835 ;
        RECT  1.485 0.925 1.890 1.085 ;
        RECT  1.225 0.805 1.485 1.085 ;
        RECT  0.785 0.925 1.225 1.085 ;
        RECT  0.640 0.925 0.785 2.500 ;
        RECT  0.625 0.925 0.640 2.940 ;
        RECT  0.385 0.925 0.625 1.085 ;
        RECT  0.380 2.340 0.625 2.940 ;
        RECT  0.125 0.820 0.385 1.085 ;
    END
END OR3X2

MACRO OR3X1
    CLASS CORE ;
    FOREIGN OR3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.630 1.105 2.635 2.290 ;
        RECT  2.370 0.810 2.630 2.290 ;
        RECT  2.225 2.130 2.370 2.290 ;
        RECT  1.965 2.130 2.225 2.730 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.545 2.110 1.715 2.400 ;
        RECT  1.225 1.760 1.545 2.400 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 1.280 1.500 1.580 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.415 0.390 1.990 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 -0.250 2.760 0.250 ;
        RECT  1.820 -0.250 2.080 0.760 ;
        RECT  1.045 -0.250 1.820 0.250 ;
        RECT  0.785 -0.250 1.045 0.405 ;
        RECT  0.000 -0.250 0.785 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.685 3.440 2.760 3.940 ;
        RECT  1.425 2.755 1.685 3.940 ;
        RECT  0.000 3.440 1.425 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.005 1.635 2.105 1.895 ;
        RECT  1.845 0.940 2.005 1.895 ;
        RECT  1.485 0.940 1.845 1.100 ;
        RECT  1.225 0.840 1.485 1.100 ;
        RECT  0.765 0.940 1.225 1.100 ;
        RECT  0.605 0.940 0.765 2.330 ;
        RECT  0.385 0.940 0.605 1.120 ;
        RECT  0.525 2.170 0.605 2.330 ;
        RECT  0.265 2.170 0.525 2.430 ;
        RECT  0.125 0.860 0.385 1.120 ;
    END
END OR3X1

MACRO OR3XL
    CLASS CORE ;
    FOREIGN OR3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.375 0.860 2.635 2.455 ;
        RECT  2.245 2.295 2.375 2.455 ;
        RECT  1.985 2.295 2.245 2.555 ;
        END
        ANTENNADIFFAREA     0.2232 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.050 1.715 2.400 ;
        RECT  1.485 2.050 1.505 2.210 ;
        RECT  1.225 1.880 1.485 2.210 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.365 1.425 1.655 ;
        RECT  1.045 1.290 1.255 1.655 ;
        RECT  0.955 1.355 1.045 1.655 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.135 1.545 0.395 2.070 ;
        RECT  0.125 1.700 0.135 1.990 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 -0.250 2.760 0.250 ;
        RECT  1.785 -0.250 2.045 0.745 ;
        RECT  1.025 -0.250 1.785 0.250 ;
        RECT  0.765 -0.250 1.025 0.405 ;
        RECT  0.000 -0.250 0.765 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.695 3.440 2.760 3.940 ;
        RECT  1.435 2.740 1.695 3.940 ;
        RECT  0.000 3.440 1.435 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.005 1.570 2.105 1.830 ;
        RECT  1.845 0.945 2.005 1.830 ;
        RECT  1.460 0.945 1.845 1.105 ;
        RECT  1.200 0.845 1.460 1.105 ;
        RECT  0.760 0.945 1.200 1.105 ;
        RECT  0.600 0.945 0.760 2.460 ;
        RECT  0.385 0.945 0.600 1.120 ;
        RECT  0.500 2.300 0.600 2.460 ;
        RECT  0.240 2.300 0.500 2.560 ;
        RECT  0.125 0.860 0.385 1.120 ;
    END
END OR3XL

MACRO OR2X8
    CLASS CORE ;
    FOREIGN OR2X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 1.105 4.015 2.585 ;
        RECT  3.960 0.610 3.965 2.585 ;
        RECT  3.705 0.610 3.960 3.020 ;
        RECT  3.700 1.005 3.705 3.020 ;
        RECT  2.945 1.005 3.700 2.200 ;
        RECT  2.940 0.610 2.945 2.200 ;
        RECT  2.860 0.610 2.940 3.050 ;
        RECT  2.685 0.610 2.860 1.295 ;
        RECT  2.680 2.035 2.860 3.050 ;
        END
        ANTENNADIFFAREA     1.5276 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.995 1.530 2.155 2.360 ;
        RECT  0.795 2.200 1.995 2.360 ;
        RECT  0.695 1.925 0.795 2.400 ;
        RECT  0.585 1.565 0.695 2.400 ;
        RECT  0.435 1.565 0.585 2.360 ;
        END
        ANTENNAGATEAREA     0.4888 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.580 1.715 1.990 ;
        RECT  1.245 1.580 1.505 1.900 ;
        END
        ANTENNAGATEAREA     0.4888 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 -0.250 4.600 0.250 ;
        RECT  4.215 -0.250 4.475 1.170 ;
        RECT  3.455 -0.250 4.215 0.250 ;
        RECT  3.195 -0.250 3.455 0.770 ;
        RECT  2.430 -0.250 3.195 0.250 ;
        RECT  2.170 -0.250 2.430 0.945 ;
        RECT  1.410 -0.250 2.170 0.250 ;
        RECT  1.150 -0.250 1.410 0.985 ;
        RECT  0.390 -0.250 1.150 0.250 ;
        RECT  0.130 -0.250 0.390 1.095 ;
        RECT  0.000 -0.250 0.130 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.470 3.440 4.600 3.940 ;
        RECT  4.210 2.080 4.470 3.940 ;
        RECT  3.450 3.440 4.210 3.940 ;
        RECT  3.190 2.420 3.450 3.940 ;
        RECT  2.405 3.440 3.190 3.940 ;
        RECT  2.145 2.950 2.405 3.940 ;
        RECT  0.730 3.440 2.145 3.940 ;
        RECT  0.470 2.610 0.730 3.940 ;
        RECT  0.000 3.440 0.470 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.495 1.540 2.640 1.800 ;
        RECT  2.335 1.190 2.495 2.745 ;
        RECT  1.920 1.190 2.335 1.350 ;
        RECT  1.555 2.585 2.335 2.745 ;
        RECT  1.660 0.825 1.920 1.350 ;
        RECT  0.900 1.190 1.660 1.350 ;
        RECT  1.295 2.585 1.555 3.185 ;
        RECT  0.740 0.835 0.900 1.350 ;
        RECT  0.640 0.835 0.740 1.095 ;
    END
END OR2X8

MACRO OR2X6
    CLASS CORE ;
    FOREIGN OR2X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 1.105 4.015 2.745 ;
        RECT  3.915 0.635 3.965 2.745 ;
        RECT  3.705 0.635 3.915 3.120 ;
        RECT  3.655 1.000 3.705 3.120 ;
        RECT  3.530 1.000 3.655 2.400 ;
        RECT  3.345 1.000 3.530 2.360 ;
        RECT  2.945 1.000 3.345 1.365 ;
        RECT  2.895 1.995 3.345 2.360 ;
        RECT  2.685 0.635 2.945 1.365 ;
        RECT  2.635 1.995 2.895 3.120 ;
        END
        ANTENNADIFFAREA     1.5776 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.005 1.635 2.070 1.895 ;
        RECT  1.845 1.635 2.005 2.360 ;
        RECT  1.810 1.635 1.845 1.895 ;
        RECT  0.795 2.200 1.845 2.360 ;
        RECT  0.665 1.925 0.795 2.400 ;
        RECT  0.585 1.695 0.665 2.400 ;
        RECT  0.455 1.695 0.585 2.360 ;
        RECT  0.405 1.695 0.455 1.955 ;
        END
        ANTENNAGATEAREA     0.3796 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.580 1.475 1.810 ;
        RECT  1.045 1.580 1.255 1.990 ;
        RECT  1.005 1.580 1.045 1.810 ;
        END
        ANTENNAGATEAREA     0.3796 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 -0.250 4.140 0.250 ;
        RECT  3.195 -0.250 3.455 0.735 ;
        RECT  2.435 -0.250 3.195 0.250 ;
        RECT  2.175 -0.250 2.435 1.000 ;
        RECT  1.415 -0.250 2.175 0.250 ;
        RECT  1.155 -0.250 1.415 1.005 ;
        RECT  0.395 -0.250 1.155 0.250 ;
        RECT  0.135 -0.250 0.395 1.075 ;
        RECT  0.000 -0.250 0.135 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 3.440 4.140 3.940 ;
        RECT  3.145 2.610 3.405 3.940 ;
        RECT  2.325 3.440 3.145 3.940 ;
        RECT  2.065 2.900 2.325 3.940 ;
        RECT  0.495 3.440 2.065 3.940 ;
        RECT  0.235 2.630 0.495 3.940 ;
        RECT  0.000 3.440 0.235 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.425 1.605 2.810 1.765 ;
        RECT  2.265 1.215 2.425 2.710 ;
        RECT  1.925 1.215 2.265 1.375 ;
        RECT  1.385 2.550 2.265 2.710 ;
        RECT  1.665 0.840 1.925 1.375 ;
        RECT  0.905 1.215 1.665 1.375 ;
        RECT  1.125 2.550 1.385 2.870 ;
        RECT  0.745 0.840 0.905 1.375 ;
        RECT  0.645 0.840 0.745 1.100 ;
    END
END OR2X6

MACRO OR2X4
    CLASS CORE ;
    FOREIGN OR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 1.080 2.205 2.290 ;
        RECT  1.990 0.620 2.035 2.290 ;
        RECT  1.965 0.620 1.990 2.400 ;
        RECT  1.775 0.620 1.965 1.320 ;
        RECT  1.865 2.050 1.965 2.400 ;
        RECT  1.605 2.050 1.865 2.990 ;
        END
        ANTENNADIFFAREA     0.7587 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.770 1.440 1.055 1.990 ;
        RECT  0.585 1.700 0.770 1.990 ;
        END
        ANTENNAGATEAREA     0.2314 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.840 ;
        RECT  0.125 1.290 0.335 1.840 ;
        RECT  0.115 1.390 0.125 1.840 ;
        END
        ANTENNAGATEAREA     0.2314 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 -0.250 2.760 0.250 ;
        RECT  2.285 -0.250 2.545 0.885 ;
        RECT  1.480 -0.250 2.285 0.250 ;
        RECT  1.220 -0.250 1.480 0.820 ;
        RECT  0.425 -0.250 1.220 0.250 ;
        RECT  0.165 -0.250 0.425 1.050 ;
        RECT  0.000 -0.250 0.165 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.375 3.440 2.760 3.940 ;
        RECT  2.115 2.585 2.375 3.940 ;
        RECT  1.315 3.440 2.115 3.940 ;
        RECT  1.055 2.550 1.315 3.940 ;
        RECT  0.000 3.440 1.055 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.415 1.560 1.695 1.820 ;
        RECT  1.255 1.050 1.415 2.350 ;
        RECT  0.935 1.050 1.255 1.210 ;
        RECT  0.425 2.190 1.255 2.350 ;
        RECT  0.675 0.885 0.935 1.210 ;
        RECT  0.165 2.080 0.425 3.020 ;
    END
END OR2X4

MACRO OR2X2
    CLASS CORE ;
    FOREIGN OR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.005 1.105 2.175 2.400 ;
        RECT  1.895 0.670 2.005 2.400 ;
        RECT  1.845 0.670 1.895 3.195 ;
        RECT  1.745 0.670 1.845 1.270 ;
        RECT  1.635 2.090 1.845 3.195 ;
        END
        ANTENNADIFFAREA     0.7004 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 1.105 1.635 ;
        END
        ANTENNAGATEAREA     0.1248 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.465 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1248 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.455 -0.250 2.300 0.250 ;
        RECT  1.195 -0.250 1.455 0.745 ;
        RECT  0.395 -0.250 1.195 0.250 ;
        RECT  0.135 -0.250 0.395 1.125 ;
        RECT  0.000 -0.250 0.135 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.345 3.440 2.300 3.940 ;
        RECT  1.085 2.440 1.345 3.940 ;
        RECT  0.000 3.440 1.085 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.455 1.580 1.655 1.840 ;
        RECT  1.295 0.950 1.455 2.260 ;
        RECT  0.905 0.950 1.295 1.110 ;
        RECT  0.745 2.100 1.295 2.260 ;
        RECT  0.645 0.850 0.905 1.110 ;
        RECT  0.585 2.100 0.745 2.425 ;
        RECT  0.415 2.265 0.585 2.425 ;
        RECT  0.155 2.265 0.415 2.865 ;
    END
END OR2X2

MACRO OR2X1
    CLASS CORE ;
    FOREIGN OR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 1.025 1.715 2.765 ;
        RECT  1.530 1.025 1.555 1.355 ;
        RECT  1.505 2.110 1.555 2.765 ;
        RECT  1.455 1.025 1.530 1.285 ;
        RECT  1.455 2.165 1.505 2.765 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.405 0.880 1.990 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.400 2.005 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 -0.250 1.840 0.250 ;
        RECT  0.900 -0.250 1.160 0.405 ;
        RECT  0.500 -0.250 0.900 0.250 ;
        RECT  0.240 -0.250 0.500 0.405 ;
        RECT  0.000 -0.250 0.240 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 3.440 1.840 3.940 ;
        RECT  1.055 3.285 1.315 3.940 ;
        RECT  0.000 3.440 1.055 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.235 1.620 1.365 1.880 ;
        RECT  1.075 0.910 1.235 2.345 ;
        RECT  0.640 0.910 1.075 1.070 ;
        RECT  0.385 2.185 1.075 2.345 ;
        RECT  0.380 0.810 0.640 1.070 ;
        RECT  0.125 2.185 0.385 2.445 ;
    END
END OR2X1

MACRO OR2XL
    CLASS CORE ;
    FOREIGN OR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.705 2.110 1.715 2.400 ;
        RECT  1.545 1.025 1.705 2.400 ;
        RECT  1.530 1.025 1.545 1.355 ;
        RECT  1.505 2.110 1.545 2.400 ;
        RECT  1.445 1.025 1.530 1.285 ;
        RECT  1.455 2.115 1.505 2.375 ;
        END
        ANTENNADIFFAREA     0.2232 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.395 0.880 1.990 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.350 1.675 0.400 1.935 ;
        RECT  0.335 1.310 0.350 1.935 ;
        RECT  0.125 1.290 0.335 1.935 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.150 -0.250 1.840 0.250 ;
        RECT  0.890 -0.250 1.150 0.405 ;
        RECT  0.490 -0.250 0.890 0.250 ;
        RECT  0.230 -0.250 0.490 0.405 ;
        RECT  0.000 -0.250 0.230 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 3.440 1.840 3.940 ;
        RECT  1.055 3.285 1.315 3.940 ;
        RECT  0.000 3.440 1.055 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.235 1.610 1.365 1.880 ;
        RECT  1.075 0.950 1.235 2.375 ;
        RECT  0.640 0.950 1.075 1.110 ;
        RECT  0.385 2.215 1.075 2.375 ;
        RECT  0.380 0.850 0.640 1.110 ;
        RECT  0.125 2.115 0.385 2.375 ;
    END
END OR2XL

MACRO NOR4BBX4
    CLASS CORE ;
    FOREIGN NOR4BBX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.430 0.880 9.535 3.030 ;
        RECT  9.190 0.590 9.430 3.030 ;
        RECT  7.050 0.590 9.190 0.825 ;
        RECT  7.050 2.830 9.190 3.030 ;
        RECT  6.670 0.535 7.050 0.825 ;
        RECT  6.290 2.830 7.050 3.090 ;
        RECT  5.850 0.585 6.670 0.825 ;
        RECT  2.680 2.830 6.290 3.030 ;
        RECT  5.590 0.535 5.850 0.825 ;
        RECT  4.770 0.585 5.590 0.825 ;
        RECT  4.510 0.535 4.770 0.825 ;
        RECT  3.690 0.585 4.510 0.825 ;
        RECT  3.430 0.535 3.690 0.825 ;
        RECT  2.610 0.585 3.430 0.825 ;
        RECT  2.420 2.595 2.680 3.195 ;
        RECT  2.350 0.550 2.610 0.825 ;
        RECT  1.530 0.595 2.350 0.825 ;
        RECT  1.270 0.550 1.530 0.825 ;
        END
        ANTENNADIFFAREA     2.4568 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.125 1.925 8.155 2.175 ;
        RECT  7.965 1.785 8.125 2.620 ;
        RECT  7.945 1.925 7.965 2.620 ;
        RECT  4.650 2.460 7.945 2.620 ;
        RECT  4.490 2.100 4.650 2.620 ;
        RECT  4.450 2.100 4.490 2.400 ;
        RECT  4.390 2.100 4.450 2.385 ;
        RECT  1.255 2.225 4.390 2.385 ;
        RECT  1.095 1.700 1.255 2.385 ;
        RECT  1.045 1.700 1.095 2.175 ;
        RECT  0.955 1.820 1.045 2.080 ;
        END
        ANTENNAGATEAREA     0.7280 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.765 1.355 7.865 1.515 ;
        RECT  7.605 1.355 7.765 2.280 ;
        RECT  5.565 2.120 7.605 2.280 ;
        RECT  5.405 1.760 5.565 2.280 ;
        RECT  3.740 1.760 5.405 1.920 ;
        RECT  3.480 1.760 3.740 2.045 ;
        RECT  1.715 1.885 3.480 2.045 ;
        RECT  1.505 1.465 1.715 2.045 ;
        RECT  1.440 1.465 1.505 1.725 ;
        END
        ANTENNAGATEAREA     0.7280 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 1.455 8.615 2.050 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.535 0.430 1.985 ;
        RECT  0.195 1.535 0.335 1.990 ;
        RECT  0.125 1.700 0.195 1.990 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.840 -0.250 9.660 0.250 ;
        RECT  7.580 -0.250 7.840 0.405 ;
        RECT  6.390 -0.250 7.580 0.250 ;
        RECT  6.130 -0.250 6.390 0.405 ;
        RECT  5.310 -0.250 6.130 0.250 ;
        RECT  5.050 -0.250 5.310 0.405 ;
        RECT  4.230 -0.250 5.050 0.250 ;
        RECT  3.970 -0.250 4.230 0.405 ;
        RECT  3.150 -0.250 3.970 0.250 ;
        RECT  2.890 -0.250 3.150 0.405 ;
        RECT  2.070 -0.250 2.890 0.250 ;
        RECT  1.810 -0.250 2.070 0.405 ;
        RECT  0.990 -0.250 1.810 0.250 ;
        RECT  0.730 -0.250 0.990 0.820 ;
        RECT  0.000 -0.250 0.730 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.375 3.440 9.660 3.940 ;
        RECT  8.115 3.285 8.375 3.940 ;
        RECT  4.815 3.440 8.115 3.940 ;
        RECT  4.215 3.285 4.815 3.940 ;
        RECT  1.020 3.440 4.215 3.940 ;
        RECT  0.760 2.890 1.020 3.940 ;
        RECT  0.000 3.440 0.760 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.795 1.115 8.955 2.525 ;
        RECT  8.645 1.115 8.795 1.275 ;
        RECT  8.685 2.265 8.795 2.525 ;
        RECT  8.385 1.015 8.645 1.275 ;
        RECT  7.385 1.015 8.385 1.175 ;
        RECT  7.285 1.015 7.385 1.720 ;
        RECT  7.225 1.015 7.285 1.915 ;
        RECT  7.125 1.460 7.225 1.915 ;
        RECT  6.385 1.755 7.125 1.915 ;
        RECT  6.805 1.415 6.905 1.575 ;
        RECT  6.645 1.035 6.805 1.575 ;
        RECT  2.780 1.035 6.645 1.195 ;
        RECT  6.225 1.415 6.385 1.915 ;
        RECT  6.125 1.415 6.225 1.735 ;
        RECT  3.260 1.415 6.125 1.575 ;
        RECT  3.000 1.415 3.260 1.675 ;
        RECT  2.270 1.485 3.000 1.645 ;
        RECT  2.520 1.035 2.780 1.305 ;
        RECT  0.770 1.035 2.520 1.195 ;
        RECT  2.010 1.375 2.270 1.645 ;
        RECT  0.610 1.035 0.770 2.335 ;
        RECT  0.385 1.035 0.610 1.195 ;
        RECT  0.395 2.175 0.610 2.335 ;
        RECT  0.135 2.175 0.395 3.115 ;
        RECT  0.125 0.595 0.385 1.195 ;
    END
END NOR4BBX4

MACRO NOR4BBX2
    CLASS CORE ;
    FOREIGN NOR4BBX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.135 0.885 6.295 2.695 ;
        RECT  5.855 0.885 6.135 1.045 ;
        RECT  5.340 2.535 6.135 2.695 ;
        RECT  5.685 0.615 5.855 1.045 ;
        RECT  3.545 0.615 5.685 0.775 ;
        RECT  5.180 2.405 5.340 2.695 ;
        RECT  4.015 2.405 5.180 2.565 ;
        RECT  3.805 2.405 4.015 2.810 ;
        RECT  3.555 2.405 3.805 2.565 ;
        RECT  3.285 2.405 3.555 3.005 ;
        RECT  3.285 0.515 3.545 0.775 ;
        RECT  2.465 0.615 3.285 0.775 ;
        RECT  2.205 0.515 2.465 0.775 ;
        END
        ANTENNADIFFAREA     1.0526 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.555 1.635 4.815 1.875 ;
        RECT  2.635 1.715 4.555 1.875 ;
        RECT  2.610 1.700 2.635 1.990 ;
        RECT  2.425 1.635 2.610 1.990 ;
        RECT  1.795 1.635 2.425 1.795 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 2.510 1.715 2.810 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.635 0.865 1.990 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.635 1.515 1.990 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.295 -0.250 6.440 0.250 ;
        RECT  6.035 -0.250 6.295 0.405 ;
        RECT  5.385 -0.250 6.035 0.250 ;
        RECT  5.125 -0.250 5.385 0.405 ;
        RECT  4.160 -0.250 5.125 0.250 ;
        RECT  3.900 -0.250 4.160 0.405 ;
        RECT  3.005 -0.250 3.900 0.250 ;
        RECT  2.745 -0.250 3.005 0.405 ;
        RECT  1.955 -0.250 2.745 0.250 ;
        RECT  1.695 -0.250 1.955 0.770 ;
        RECT  0.935 -0.250 1.695 0.250 ;
        RECT  0.675 -0.250 0.935 1.095 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.985 3.440 6.440 3.940 ;
        RECT  4.725 2.745 4.985 3.940 ;
        RECT  2.055 3.440 4.725 3.940 ;
        RECT  1.895 2.560 2.055 3.940 ;
        RECT  0.895 3.440 1.895 3.940 ;
        RECT  0.635 2.170 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.795 1.225 5.955 2.305 ;
        RECT  5.500 1.225 5.795 1.385 ;
        RECT  2.975 2.055 5.795 2.215 ;
        RECT  5.455 1.565 5.615 1.825 ;
        RECT  5.340 0.955 5.500 1.385 ;
        RECT  5.155 1.565 5.455 1.725 ;
        RECT  3.715 0.955 5.340 1.115 ;
        RECT  4.995 1.295 5.155 1.725 ;
        RECT  4.195 1.295 4.995 1.455 ;
        RECT  3.935 1.295 4.195 1.535 ;
        RECT  3.205 1.375 3.935 1.535 ;
        RECT  3.455 0.955 3.715 1.195 ;
        RECT  1.445 0.955 3.455 1.115 ;
        RECT  3.155 1.300 3.205 1.535 ;
        RECT  2.945 1.295 3.155 1.535 ;
        RECT  2.815 2.055 2.975 2.330 ;
        RECT  0.285 1.295 2.945 1.455 ;
        RECT  1.145 2.170 2.815 2.330 ;
        RECT  1.185 0.855 1.445 1.115 ;
        RECT  0.285 0.835 0.425 1.095 ;
        RECT  0.285 2.170 0.385 2.770 ;
        RECT  0.125 0.835 0.285 2.770 ;
    END
END NOR4BBX2

MACRO NOR4BBX1
    CLASS CORE ;
    FOREIGN NOR4BBX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 0.695 3.565 2.930 ;
        RECT  2.320 0.695 3.405 0.855 ;
        RECT  2.635 2.770 3.405 2.930 ;
        RECT  2.600 2.770 2.635 3.220 ;
        RECT  2.425 2.675 2.600 3.220 ;
        RECT  2.340 2.675 2.425 2.995 ;
        RECT  2.060 0.640 2.320 0.925 ;
        RECT  1.370 0.765 2.060 0.925 ;
        RECT  1.110 0.765 1.370 1.035 ;
        END
        ANTENNADIFFAREA     0.7120 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.155 1.700 1.255 1.990 ;
        RECT  1.045 1.410 1.155 1.990 ;
        RECT  0.910 1.410 1.045 1.865 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.265 1.715 1.795 ;
        RECT  1.365 1.265 1.505 1.525 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.650 3.225 2.100 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.290 0.385 1.795 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.920 -0.250 3.680 0.250 ;
        RECT  2.660 -0.250 2.920 0.405 ;
        RECT  1.770 -0.250 2.660 0.250 ;
        RECT  1.510 -0.250 1.770 0.405 ;
        RECT  0.820 -0.250 1.510 0.250 ;
        RECT  0.560 -0.250 0.820 0.405 ;
        RECT  0.000 -0.250 0.560 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.365 3.440 3.680 3.940 ;
        RECT  3.105 3.285 3.365 3.940 ;
        RECT  1.105 3.440 3.105 3.940 ;
        RECT  0.845 2.540 1.105 3.940 ;
        RECT  0.000 3.440 0.845 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.950 2.310 3.210 2.570 ;
        RECT  3.040 1.035 3.200 1.365 ;
        RECT  2.705 1.205 3.040 1.365 ;
        RECT  2.705 2.310 2.950 2.470 ;
        RECT  2.545 1.205 2.705 2.470 ;
        RECT  2.155 1.205 2.545 1.365 ;
        RECT  2.205 1.585 2.365 2.335 ;
        RECT  0.730 2.175 2.205 2.335 ;
        RECT  1.895 1.105 2.155 1.365 ;
        RECT  0.570 0.950 0.730 2.335 ;
        RECT  0.385 0.950 0.570 1.110 ;
        RECT  0.125 2.035 0.570 2.335 ;
        RECT  0.125 0.850 0.385 1.110 ;
    END
END NOR4BBX1

MACRO NOR4BBXL
    CLASS CORE ;
    FOREIGN NOR4BBXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.530 1.700 3.555 1.990 ;
        RECT  3.520 0.695 3.530 1.990 ;
        RECT  3.370 0.695 3.520 2.735 ;
        RECT  2.500 0.695 3.370 0.855 ;
        RECT  3.360 1.700 3.370 2.735 ;
        RECT  3.345 1.700 3.360 1.990 ;
        RECT  2.370 2.575 3.360 2.735 ;
        RECT  2.240 0.695 2.500 1.025 ;
        RECT  1.400 0.865 2.240 1.025 ;
        RECT  1.140 0.865 1.400 1.125 ;
        END
        ANTENNADIFFAREA     0.5781 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.700 1.255 1.990 ;
        RECT  1.045 1.470 1.180 1.990 ;
        RECT  0.935 1.470 1.045 1.965 ;
        END
        ANTENNAGATEAREA     0.1131 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.290 1.715 1.780 ;
        RECT  1.415 1.305 1.505 1.565 ;
        END
        ANTENNAGATEAREA     0.1131 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.570 3.145 2.050 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.290 0.385 1.805 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 -0.250 3.680 0.250 ;
        RECT  2.980 -0.250 3.240 0.405 ;
        RECT  1.640 -0.250 2.980 0.250 ;
        RECT  1.380 -0.250 1.640 0.405 ;
        RECT  0.820 -0.250 1.380 0.250 ;
        RECT  0.560 -0.250 0.820 0.405 ;
        RECT  0.000 -0.250 0.560 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.140 3.440 3.680 3.940 ;
        RECT  2.880 3.285 3.140 3.940 ;
        RECT  1.105 3.440 2.880 3.940 ;
        RECT  0.845 2.550 1.105 3.940 ;
        RECT  0.000 3.440 0.845 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.030 1.035 3.190 1.385 ;
        RECT  2.705 2.235 3.180 2.395 ;
        RECT  2.705 1.225 3.030 1.385 ;
        RECT  2.545 1.225 2.705 2.395 ;
        RECT  2.055 1.225 2.545 1.415 ;
        RECT  2.205 1.715 2.365 1.975 ;
        RECT  2.145 1.815 2.205 1.975 ;
        RECT  1.985 1.815 2.145 2.335 ;
        RECT  1.895 1.225 2.055 1.495 ;
        RECT  0.755 2.175 1.985 2.335 ;
        RECT  0.595 0.950 0.755 2.335 ;
        RECT  0.385 0.950 0.595 1.110 ;
        RECT  0.385 2.175 0.595 2.335 ;
        RECT  0.125 0.850 0.385 1.110 ;
        RECT  0.125 2.140 0.385 2.400 ;
    END
END NOR4BBXL

MACRO NOR4BX4
    CLASS CORE ;
    FOREIGN NOR4BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.365 0.585 8.615 3.100 ;
        RECT  6.930 0.585 8.365 0.825 ;
        RECT  7.050 2.860 8.365 3.100 ;
        RECT  6.645 2.860 7.050 3.150 ;
        RECT  6.670 0.535 6.930 0.825 ;
        RECT  5.850 0.585 6.670 0.825 ;
        RECT  2.910 2.860 6.645 3.100 ;
        RECT  5.590 0.535 5.850 0.825 ;
        RECT  4.770 0.585 5.590 0.825 ;
        RECT  4.510 0.535 4.770 0.825 ;
        RECT  3.690 0.585 4.510 0.825 ;
        RECT  3.430 0.535 3.690 0.825 ;
        RECT  2.610 0.585 3.430 0.825 ;
        RECT  2.520 2.860 2.910 3.140 ;
        RECT  2.350 0.535 2.610 0.825 ;
        RECT  1.530 0.585 2.350 0.825 ;
        RECT  1.270 0.535 1.530 0.825 ;
        END
        ANTENNADIFFAREA     1.8848 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.155 1.820 8.175 2.080 ;
        RECT  8.105 1.820 8.155 2.400 ;
        RECT  7.945 1.820 8.105 2.565 ;
        RECT  7.915 1.820 7.945 2.080 ;
        RECT  5.005 2.405 7.945 2.565 ;
        RECT  4.405 2.305 5.005 2.565 ;
        RECT  4.030 2.405 4.405 2.565 ;
        RECT  3.870 2.405 4.030 2.675 ;
        RECT  1.325 2.515 3.870 2.675 ;
        RECT  1.165 1.585 1.325 2.675 ;
        RECT  1.065 1.585 1.165 1.845 ;
        END
        ANTENNAGATEAREA     0.7280 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.920 1.275 8.180 1.535 ;
        RECT  7.725 1.375 7.920 1.535 ;
        RECT  7.565 1.375 7.725 2.105 ;
        RECT  5.945 1.945 7.565 2.105 ;
        RECT  5.685 1.760 5.945 2.105 ;
        RECT  3.740 1.760 5.685 1.920 ;
        RECT  3.690 1.760 3.740 2.045 ;
        RECT  3.480 1.760 3.690 2.335 ;
        RECT  1.770 2.170 3.480 2.335 ;
        RECT  1.610 1.445 1.770 2.335 ;
        RECT  1.505 1.445 1.610 1.990 ;
        END
        ANTENNAGATEAREA     0.7280 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.125 1.415 7.385 1.700 ;
        RECT  6.500 1.415 7.125 1.575 ;
        RECT  6.240 1.415 6.500 1.700 ;
        RECT  3.260 1.415 6.240 1.575 ;
        RECT  3.000 1.415 3.260 1.675 ;
        RECT  2.300 1.515 3.000 1.675 ;
        RECT  2.175 1.445 2.300 1.925 ;
        RECT  2.040 1.445 2.175 1.990 ;
        RECT  1.965 1.700 2.040 1.990 ;
        END
        ANTENNAGATEAREA     0.7280 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.580 0.545 1.990 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.470 -0.250 8.740 0.250 ;
        RECT  7.210 -0.250 7.470 0.405 ;
        RECT  6.390 -0.250 7.210 0.250 ;
        RECT  6.130 -0.250 6.390 0.405 ;
        RECT  5.310 -0.250 6.130 0.250 ;
        RECT  5.050 -0.250 5.310 0.405 ;
        RECT  4.230 -0.250 5.050 0.250 ;
        RECT  3.970 -0.250 4.230 0.405 ;
        RECT  3.150 -0.250 3.970 0.250 ;
        RECT  2.890 -0.250 3.150 0.405 ;
        RECT  2.070 -0.250 2.890 0.250 ;
        RECT  1.810 -0.250 2.070 0.405 ;
        RECT  0.990 -0.250 1.810 0.250 ;
        RECT  0.730 -0.250 0.990 0.820 ;
        RECT  0.000 -0.250 0.730 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.375 3.440 8.740 3.940 ;
        RECT  8.115 3.285 8.375 3.940 ;
        RECT  4.445 3.440 8.115 3.940 ;
        RECT  4.185 3.285 4.445 3.940 ;
        RECT  1.260 3.440 4.185 3.940 ;
        RECT  1.000 2.955 1.260 3.940 ;
        RECT  0.000 3.440 1.000 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.780 1.005 7.700 1.165 ;
        RECT  2.520 1.005 2.780 1.310 ;
        RECT  0.885 1.005 2.520 1.165 ;
        RECT  0.725 1.005 0.885 2.390 ;
        RECT  0.450 1.005 0.725 1.165 ;
        RECT  0.675 2.225 0.725 2.390 ;
        RECT  0.415 2.225 0.675 3.165 ;
        RECT  0.190 0.565 0.450 1.165 ;
    END
END NOR4BX4

MACRO NOR4BX2
    CLASS CORE ;
    FOREIGN NOR4BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 0.980 4.935 2.810 ;
        RECT  4.775 0.980 4.885 3.040 ;
        RECT  4.305 0.980 4.775 1.140 ;
        RECT  4.725 2.335 4.775 3.040 ;
        RECT  2.575 2.880 4.725 3.040 ;
        RECT  3.990 0.875 4.305 1.140 ;
        RECT  3.355 0.875 3.990 1.035 ;
        RECT  3.255 0.775 3.355 1.035 ;
        RECT  3.095 0.635 3.255 1.035 ;
        RECT  2.415 0.635 3.095 0.795 ;
        RECT  2.315 2.880 2.575 3.140 ;
        RECT  2.150 0.535 2.415 0.795 ;
        RECT  1.335 0.635 2.150 0.795 ;
        RECT  1.075 0.535 1.335 0.795 ;
        END
        ANTENNADIFFAREA     1.1874 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.635 4.115 1.895 ;
        RECT  3.965 1.635 4.015 1.990 ;
        RECT  3.855 1.635 3.965 2.330 ;
        RECT  3.805 1.685 3.855 2.330 ;
        RECT  1.050 2.170 3.805 2.330 ;
        RECT  0.890 1.635 1.050 2.330 ;
        END
        ANTENNAGATEAREA     0.4264 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.325 3.570 1.585 ;
        RECT  3.310 1.325 3.555 1.990 ;
        RECT  3.305 1.375 3.310 1.990 ;
        RECT  1.580 1.830 3.305 1.990 ;
        RECT  1.420 1.325 1.580 1.990 ;
        RECT  1.320 1.325 1.420 1.585 ;
        END
        ANTENNAGATEAREA     0.4264 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.290 3.095 1.625 ;
        RECT  2.830 1.325 2.885 1.625 ;
        RECT  2.060 1.465 2.830 1.625 ;
        RECT  1.800 1.325 2.060 1.625 ;
        END
        ANTENNAGATEAREA     0.4264 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.105 1.275 0.335 1.810 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.855 -0.250 5.060 0.250 ;
        RECT  4.595 -0.250 4.855 0.800 ;
        RECT  3.905 -0.250 4.595 0.250 ;
        RECT  3.645 -0.250 3.905 0.405 ;
        RECT  2.965 -0.250 3.645 0.250 ;
        RECT  2.705 -0.250 2.965 0.405 ;
        RECT  1.875 -0.250 2.705 0.250 ;
        RECT  1.615 -0.250 1.875 0.405 ;
        RECT  0.785 -0.250 1.615 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.090 3.440 5.060 3.940 ;
        RECT  3.830 3.285 4.090 3.940 ;
        RECT  1.070 3.440 3.830 3.940 ;
        RECT  0.810 2.880 1.070 3.940 ;
        RECT  0.000 3.440 0.810 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.545 1.320 4.595 1.580 ;
        RECT  4.385 1.320 4.545 2.670 ;
        RECT  4.335 1.320 4.385 1.580 ;
        RECT  0.385 2.510 4.385 2.670 ;
        RECT  2.325 0.985 2.585 1.285 ;
        RECT  0.675 0.985 2.325 1.145 ;
        RECT  0.515 0.835 0.675 2.160 ;
        RECT  0.125 0.835 0.515 1.095 ;
        RECT  0.385 2.000 0.515 2.160 ;
        RECT  0.125 2.000 0.385 2.685 ;
    END
END NOR4BX2

MACRO NOR4BX1
    CLASS CORE ;
    FOREIGN NOR4BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 0.920 3.095 2.585 ;
        RECT  2.450 0.920 2.815 1.080 ;
        RECT  2.555 2.420 2.815 2.585 ;
        RECT  2.295 2.420 2.555 3.020 ;
        RECT  2.055 0.820 2.450 1.080 ;
        RECT  1.530 0.920 2.055 1.080 ;
        RECT  1.105 0.820 1.530 1.080 ;
        END
        ANTENNADIFFAREA     0.7125 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.115 1.700 1.255 1.990 ;
        RECT  0.855 1.475 1.115 1.990 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 1.360 1.715 1.990 ;
        RECT  1.335 1.360 1.435 1.520 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 1.290 2.175 1.750 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.380 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.865 -0.250 3.220 0.250 ;
        RECT  2.605 -0.250 2.865 0.405 ;
        RECT  1.765 -0.250 2.605 0.250 ;
        RECT  1.505 -0.250 1.765 0.405 ;
        RECT  0.815 -0.250 1.505 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.115 3.440 3.220 3.940 ;
        RECT  0.855 2.615 1.115 3.940 ;
        RECT  0.000 3.440 0.855 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.535 1.655 2.635 1.915 ;
        RECT  2.375 1.655 2.535 2.235 ;
        RECT  2.055 2.075 2.375 2.235 ;
        RECT  1.895 2.075 2.055 2.435 ;
        RECT  0.675 2.275 1.895 2.435 ;
        RECT  0.515 1.040 0.675 2.435 ;
        RECT  0.385 1.040 0.515 1.200 ;
        RECT  0.385 2.220 0.515 2.435 ;
        RECT  0.125 0.940 0.385 1.200 ;
        RECT  0.125 2.220 0.385 2.480 ;
    END
END NOR4BX1

MACRO NOR4BXL
    CLASS CORE ;
    FOREIGN NOR4BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.040 1.290 3.095 2.465 ;
        RECT  2.880 0.945 3.040 2.465 ;
        RECT  2.520 0.945 2.880 1.105 ;
        RECT  2.560 2.305 2.880 2.465 ;
        RECT  2.300 2.305 2.560 2.565 ;
        RECT  2.450 0.845 2.520 1.105 ;
        RECT  2.260 0.705 2.450 1.105 ;
        RECT  1.400 0.705 2.260 0.865 ;
        RECT  1.140 0.605 1.400 0.865 ;
        END
        ANTENNADIFFAREA     0.4681 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.010 1.550 1.270 2.020 ;
        END
        ANTENNAGATEAREA     0.1131 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.665 1.290 1.715 1.580 ;
        RECT  1.515 1.120 1.665 1.580 ;
        RECT  1.505 1.070 1.515 1.580 ;
        RECT  1.255 1.070 1.505 1.330 ;
        END
        ANTENNAGATEAREA     0.1131 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.170 1.290 2.175 1.580 ;
        RECT  2.055 1.290 2.170 1.740 ;
        RECT  1.895 1.265 2.055 1.740 ;
        END
        ANTENNAGATEAREA     0.1131 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.380 1.480 0.410 1.740 ;
        RECT  0.130 1.230 0.380 1.740 ;
        RECT  0.125 1.290 0.130 1.580 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.220 0.250 ;
        RECT  2.835 -0.250 3.095 0.765 ;
        RECT  1.980 -0.250 2.835 0.250 ;
        RECT  1.720 -0.250 1.980 0.405 ;
        RECT  0.790 -0.250 1.720 0.250 ;
        RECT  0.170 -0.250 0.790 0.405 ;
        RECT  0.000 -0.250 0.170 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.090 3.440 3.220 3.940 ;
        RECT  0.830 2.555 1.090 3.940 ;
        RECT  0.000 3.440 0.830 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.530 1.385 2.630 1.645 ;
        RECT  2.370 1.385 2.530 2.120 ;
        RECT  1.920 1.960 2.370 2.120 ;
        RECT  1.760 1.960 1.920 2.360 ;
        RECT  0.750 2.200 1.760 2.360 ;
        RECT  0.750 1.035 0.830 1.295 ;
        RECT  0.590 1.035 0.750 2.360 ;
        RECT  0.570 1.035 0.590 1.295 ;
        RECT  0.180 1.955 0.590 2.215 ;
    END
END NOR4BXL

MACRO NOR3BX4
    CLASS CORE ;
    FOREIGN NOR3BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.755 2.515 4.015 3.145 ;
        RECT  3.705 0.640 3.965 0.900 ;
        RECT  1.755 2.515 3.755 2.755 ;
        RECT  2.885 0.660 3.705 0.900 ;
        RECT  2.625 0.640 2.885 0.900 ;
        RECT  1.805 0.660 2.625 0.900 ;
        RECT  1.545 0.640 1.805 0.900 ;
        RECT  1.495 2.515 1.755 3.145 ;
        RECT  0.365 0.660 1.545 0.900 ;
        RECT  0.365 2.515 1.495 2.755 ;
        RECT  0.125 0.660 0.365 2.755 ;
        END
        ANTENNADIFFAREA     1.7969 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 1.775 4.985 2.035 ;
        RECT  4.725 1.775 4.935 2.335 ;
        RECT  2.930 2.175 4.725 2.335 ;
        RECT  2.770 1.775 2.930 2.335 ;
        RECT  0.795 2.175 2.770 2.335 ;
        RECT  0.610 1.700 0.795 2.335 ;
        RECT  0.585 1.700 0.610 2.035 ;
        END
        ANTENNAGATEAREA     0.7852 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 0.950 4.735 1.240 ;
        RECT  4.265 0.880 4.475 1.240 ;
        RECT  3.710 1.080 4.265 1.240 ;
        RECT  3.450 1.080 3.710 1.630 ;
        RECT  2.220 1.080 3.450 1.240 ;
        RECT  1.960 1.080 2.220 1.630 ;
        RECT  0.895 1.080 1.960 1.240 ;
        RECT  0.735 1.080 0.895 1.520 ;
        RECT  0.635 1.260 0.735 1.520 ;
        END
        ANTENNAGATEAREA     0.7852 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.865 1.485 6.315 1.990 ;
        END
        ANTENNAGATEAREA     0.3016 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.295 -0.250 6.440 0.250 ;
        RECT  6.035 -0.250 6.295 1.055 ;
        RECT  5.245 -0.250 6.035 0.250 ;
        RECT  4.985 -0.250 5.245 1.140 ;
        RECT  4.505 -0.250 4.985 0.250 ;
        RECT  4.245 -0.250 4.505 0.405 ;
        RECT  3.425 -0.250 4.245 0.250 ;
        RECT  3.165 -0.250 3.425 0.405 ;
        RECT  2.345 -0.250 3.165 0.250 ;
        RECT  2.085 -0.250 2.345 0.405 ;
        RECT  1.265 -0.250 2.085 0.250 ;
        RECT  1.005 -0.250 1.265 0.405 ;
        RECT  0.000 -0.250 1.005 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.295 3.440 6.440 3.940 ;
        RECT  6.035 2.205 6.295 3.940 ;
        RECT  5.195 3.440 6.035 3.940 ;
        RECT  4.935 2.540 5.195 3.940 ;
        RECT  2.885 3.440 4.935 3.940 ;
        RECT  2.625 2.935 2.885 3.940 ;
        RECT  0.625 3.440 2.625 3.940 ;
        RECT  0.365 2.935 0.625 3.940 ;
        RECT  0.000 3.440 0.365 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.665 0.805 5.785 1.065 ;
        RECT  5.665 2.205 5.785 2.805 ;
        RECT  5.505 0.805 5.665 2.805 ;
        RECT  5.445 0.805 5.505 1.580 ;
        RECT  4.195 1.420 5.445 1.580 ;
        RECT  4.095 1.420 4.195 1.680 ;
        RECT  3.935 1.420 4.095 1.995 ;
        RECT  3.270 1.835 3.935 1.995 ;
        RECT  3.110 1.430 3.270 1.995 ;
        RECT  2.590 1.430 3.110 1.590 ;
        RECT  2.430 1.430 2.590 1.990 ;
        RECT  1.585 1.830 2.430 1.990 ;
        RECT  1.325 1.730 1.585 1.990 ;
    END
END NOR3BX4

MACRO NOR3BX2
    CLASS CORE ;
    FOREIGN NOR3BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.745 0.565 2.005 1.165 ;
        RECT  0.925 0.935 1.745 1.095 ;
        RECT  1.615 2.930 1.715 3.220 ;
        RECT  1.505 2.580 1.615 3.220 ;
        RECT  1.355 2.580 1.505 3.180 ;
        RECT  0.265 2.580 1.355 2.740 ;
        RECT  0.825 0.495 0.925 1.095 ;
        RECT  0.665 0.495 0.825 1.165 ;
        RECT  0.585 0.695 0.665 1.165 ;
        RECT  0.335 1.005 0.585 1.165 ;
        RECT  0.265 1.005 0.335 1.355 ;
        RECT  0.105 1.005 0.265 2.740 ;
        END
        ANTENNADIFFAREA     1.0190 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.615 1.775 2.775 2.400 ;
        RECT  0.795 2.240 2.615 2.400 ;
        RECT  0.605 2.110 0.795 2.400 ;
        RECT  0.445 1.775 0.605 2.400 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 1.405 2.095 1.665 ;
        RECT  1.255 1.405 1.935 1.565 ;
        RECT  1.135 1.290 1.255 1.580 ;
        RECT  1.045 1.290 1.135 1.680 ;
        RECT  0.875 1.405 1.045 1.680 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.295 1.450 3.555 2.025 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 -0.250 3.680 0.250 ;
        RECT  2.260 -0.250 2.520 1.140 ;
        RECT  1.465 -0.250 2.260 0.250 ;
        RECT  1.205 -0.250 1.465 0.745 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 3.440 3.680 3.940 ;
        RECT  2.510 2.595 2.770 3.940 ;
        RECT  0.455 3.440 2.510 3.940 ;
        RECT  0.195 2.945 0.455 3.940 ;
        RECT  0.000 3.440 0.195 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.215 2.205 3.475 2.805 ;
        RECT  3.115 2.205 3.215 2.365 ;
        RECT  3.060 1.355 3.115 2.365 ;
        RECT  2.955 0.985 3.060 2.365 ;
        RECT  2.800 0.985 2.955 1.515 ;
        RECT  2.435 1.355 2.800 1.515 ;
        RECT  2.275 1.355 2.435 2.035 ;
        RECT  1.615 1.875 2.275 2.035 ;
        RECT  1.355 1.775 1.615 2.035 ;
    END
END NOR3BX2

MACRO NOR3BX1
    CLASS CORE ;
    FOREIGN NOR3BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 0.880 2.635 2.695 ;
        RECT  2.425 0.880 2.475 1.355 ;
        RECT  2.450 2.335 2.475 2.695 ;
        RECT  2.425 2.335 2.450 2.810 ;
        RECT  2.375 0.955 2.425 1.215 ;
        RECT  2.290 2.535 2.425 2.810 ;
        RECT  1.530 1.055 2.375 1.215 ;
        RECT  2.030 2.535 2.290 3.135 ;
        RECT  1.965 2.745 2.030 2.995 ;
        RECT  1.270 0.955 1.530 1.215 ;
        END
        ANTENNADIFFAREA     0.6730 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.405 1.255 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.395 1.810 1.655 ;
        RECT  1.505 1.395 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.500 1.465 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 -0.250 2.760 0.250 ;
        RECT  1.820 -0.250 2.080 0.825 ;
        RECT  0.990 -0.250 1.820 0.250 ;
        RECT  0.730 -0.250 0.990 1.135 ;
        RECT  0.000 -0.250 0.730 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 3.440 2.760 3.940 ;
        RECT  0.870 2.535 1.130 3.940 ;
        RECT  0.000 3.440 0.870 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.195 1.705 2.295 1.965 ;
        RECT  2.035 1.705 2.195 2.330 ;
        RECT  0.590 2.170 2.035 2.330 ;
        RECT  0.330 2.170 0.590 2.430 ;
        RECT  0.320 1.025 0.420 1.285 ;
        RECT  0.320 2.170 0.330 2.330 ;
        RECT  0.160 1.025 0.320 2.330 ;
    END
END NOR3BX1

MACRO NOR3BXL
    CLASS CORE ;
    FOREIGN NOR3BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 0.470 2.175 2.670 ;
        RECT  1.915 0.535 1.965 0.965 ;
        RECT  1.915 2.335 1.965 2.670 ;
        RECT  1.260 0.805 1.915 0.965 ;
        RECT  1.000 0.705 1.260 0.965 ;
        END
        ANTENNADIFFAREA     0.5877 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.655 0.880 1.915 ;
        RECT  0.585 1.555 0.835 2.025 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 1.420 1.475 1.840 ;
        RECT  1.255 1.420 1.315 1.580 ;
        RECT  1.045 1.290 1.255 1.580 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.790 0.555 3.050 ;
        RECT  0.150 2.790 0.335 3.220 ;
        RECT  0.125 2.930 0.150 3.220 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.610 -0.250 2.300 0.250 ;
        RECT  0.670 -0.250 1.610 0.405 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.995 3.440 2.300 3.940 ;
        RECT  0.735 2.800 0.995 3.940 ;
        RECT  0.000 3.440 0.735 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.745 2.930 2.005 3.190 ;
        RECT  1.585 2.930 1.745 3.090 ;
        RECT  1.425 2.345 1.585 3.090 ;
        RECT  0.385 2.345 1.425 2.505 ;
        RECT  0.285 0.605 0.385 0.865 ;
        RECT  0.285 2.345 0.385 2.605 ;
        RECT  0.125 0.605 0.285 2.605 ;
    END
END NOR3BXL

MACRO NOR2BX4
    CLASS CORE ;
    FOREIGN NOR2BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.415 0.885 3.555 2.585 ;
        RECT  3.345 0.885 3.415 2.930 ;
        RECT  2.425 0.885 3.345 1.085 ;
        RECT  3.155 2.330 3.345 2.930 ;
        RECT  1.775 2.330 3.155 2.530 ;
        RECT  2.165 0.815 2.425 1.085 ;
        RECT  1.405 0.885 2.165 1.085 ;
        RECT  1.515 2.330 1.775 2.930 ;
        RECT  1.145 0.825 1.405 1.085 ;
        END
        ANTENNADIFFAREA     1.4320 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 1.630 2.635 1.790 ;
        RECT  2.325 1.630 2.485 2.120 ;
        RECT  1.305 1.960 2.325 2.120 ;
        RECT  1.145 1.625 1.305 2.120 ;
        RECT  1.045 1.625 1.145 1.990 ;
        RECT  0.865 1.625 1.045 1.785 ;
        END
        ANTENNAGATEAREA     0.6474 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.455 0.345 2.060 ;
        END
        ANTENNAGATEAREA     0.2522 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 -0.250 3.680 0.250 ;
        RECT  2.715 -0.250 2.975 0.405 ;
        RECT  1.915 -0.250 2.715 0.250 ;
        RECT  1.655 -0.250 1.915 0.685 ;
        RECT  0.895 -0.250 1.655 0.250 ;
        RECT  0.635 -0.250 0.895 0.840 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.595 3.440 3.680 3.940 ;
        RECT  2.335 2.750 2.595 3.940 ;
        RECT  0.925 3.440 2.335 3.940 ;
        RECT  0.665 2.885 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.985 1.270 3.145 1.530 ;
        RECT  1.895 1.285 2.985 1.445 ;
        RECT  1.635 1.285 1.895 1.760 ;
        RECT  0.690 1.285 1.635 1.445 ;
        RECT  0.685 1.105 0.690 1.445 ;
        RECT  0.525 1.105 0.685 2.475 ;
        RECT  0.385 1.105 0.525 1.265 ;
        RECT  0.385 2.315 0.525 2.475 ;
        RECT  0.125 0.665 0.385 1.265 ;
        RECT  0.125 2.315 0.385 2.915 ;
    END
END NOR2BX4

MACRO NOR2BX2
    CLASS CORE ;
    FOREIGN NOR2BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.580 1.515 2.635 2.335 ;
        RECT  2.420 1.060 2.580 2.505 ;
        RECT  2.085 1.060 2.420 1.220 ;
        RECT  1.715 2.345 2.420 2.505 ;
        RECT  1.825 0.620 2.085 1.220 ;
        RECT  1.505 2.345 1.715 2.810 ;
        RECT  1.380 2.345 1.505 2.605 ;
        END
        ANTENNADIFFAREA     0.6384 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 1.595 2.240 2.020 ;
        RECT  1.255 1.860 2.080 2.020 ;
        RECT  1.110 1.290 1.255 2.020 ;
        RECT  1.065 1.280 1.110 2.020 ;
        RECT  1.045 1.280 1.065 1.765 ;
        RECT  0.950 1.280 1.045 1.540 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.510 0.430 1.985 ;
        RECT  0.175 1.510 0.335 1.990 ;
        RECT  0.125 1.700 0.175 1.990 ;
        END
        ANTENNAGATEAREA     0.1248 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.595 -0.250 2.760 0.250 ;
        RECT  2.335 -0.250 2.595 0.840 ;
        RECT  1.540 -0.250 2.335 0.250 ;
        RECT  1.280 -0.250 1.540 0.755 ;
        RECT  0.000 -0.250 1.280 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.500 3.440 2.760 3.940 ;
        RECT  2.240 2.885 2.500 3.940 ;
        RECT  0.925 3.440 2.240 3.940 ;
        RECT  0.665 3.285 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.600 1.420 1.700 1.680 ;
        RECT  1.440 0.935 1.600 1.680 ;
        RECT  1.000 0.935 1.440 1.095 ;
        RECT  0.770 0.510 1.000 1.095 ;
        RECT  0.740 0.510 0.770 2.410 ;
        RECT  0.610 0.935 0.740 2.410 ;
        RECT  0.385 2.250 0.610 2.410 ;
        RECT  0.125 2.250 0.385 2.510 ;
    END
END NOR2BX2

MACRO NOR2BX1
    CLASS CORE ;
    FOREIGN NOR2BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 0.880 1.730 2.285 ;
        RECT  1.660 0.880 1.715 2.585 ;
        RECT  1.570 0.880 1.660 2.720 ;
        RECT  1.505 0.880 1.570 1.170 ;
        RECT  1.400 2.120 1.570 2.720 ;
        RECT  1.040 0.920 1.505 1.080 ;
        END
        ANTENNADIFFAREA     0.4872 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.600 0.880 2.335 ;
        RECT  0.720 1.600 0.795 2.400 ;
        RECT  0.585 1.925 0.720 2.400 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.380 1.600 0.400 1.860 ;
        RECT  0.115 1.530 0.380 1.990 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 -0.250 1.840 0.250 ;
        RECT  0.980 -0.250 1.700 0.405 ;
        RECT  0.000 -0.250 0.980 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 3.440 1.840 3.940 ;
        RECT  0.640 3.285 0.900 3.940 ;
        RECT  0.000 3.440 0.640 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.220 1.590 1.390 1.865 ;
        RECT  1.060 1.260 1.220 2.740 ;
        RECT  0.800 1.260 1.060 1.420 ;
        RECT  0.385 2.580 1.060 2.740 ;
        RECT  0.640 0.620 0.800 1.420 ;
        RECT  0.390 0.620 0.640 0.780 ;
        RECT  0.130 0.520 0.390 0.780 ;
        RECT  0.125 2.540 0.385 2.800 ;
    END
END NOR2BX1

MACRO NOR2BXL
    CLASS CORE ;
    FOREIGN NOR2BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.570 0.975 1.730 2.425 ;
        RECT  1.225 0.975 1.570 1.135 ;
        RECT  1.505 2.110 1.570 2.425 ;
        RECT  1.400 2.165 1.505 2.425 ;
        END
        ANTENNADIFFAREA     0.3765 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.660 0.875 2.335 ;
        RECT  0.715 1.660 0.795 2.400 ;
        RECT  0.585 1.925 0.715 2.400 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.340 1.660 0.395 1.920 ;
        RECT  0.125 1.660 0.340 2.205 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 -0.250 1.840 0.250 ;
        RECT  0.975 -0.250 1.235 0.405 ;
        RECT  0.000 -0.250 0.975 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 3.440 1.840 3.940 ;
        RECT  0.635 2.945 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.220 1.645 1.385 1.920 ;
        RECT  1.060 1.320 1.220 2.740 ;
        RECT  0.385 1.320 1.060 1.480 ;
        RECT  0.385 2.580 1.060 2.740 ;
        RECT  0.225 0.600 0.385 1.480 ;
        RECT  0.125 2.540 0.385 2.800 ;
        RECT  0.125 0.600 0.225 0.860 ;
    END
END NOR2BXL

MACRO NOR4X8
    CLASS CORE ;
    FOREIGN NOR4X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.100 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.665 0.585 15.975 3.105 ;
        RECT  15.305 0.585 15.665 1.580 ;
        RECT  3.425 2.705 15.665 3.105 ;
        RECT  14.560 0.585 15.305 0.885 ;
        RECT  12.700 0.585 14.560 0.865 ;
        RECT  0.925 0.585 12.700 0.885 ;
        RECT  1.850 2.815 3.425 3.105 ;
        RECT  0.665 0.585 0.925 1.110 ;
        END
        ANTENNADIFFAREA     4.0956 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.325 1.815 15.485 2.485 ;
        RECT  12.270 2.325 15.325 2.485 ;
        RECT  12.010 2.265 12.270 2.525 ;
        RECT  8.175 2.325 12.010 2.485 ;
        RECT  7.915 2.225 8.175 2.485 ;
        RECT  4.175 2.325 7.915 2.485 ;
        RECT  3.915 2.225 4.175 2.485 ;
        RECT  3.245 2.325 3.915 2.485 ;
        RECT  3.085 2.325 3.245 2.600 ;
        RECT  0.585 2.440 3.085 2.600 ;
        RECT  0.425 1.805 0.585 2.600 ;
        RECT  0.325 1.805 0.425 2.400 ;
        RECT  0.125 2.110 0.325 2.400 ;
        END
        ANTENNAGATEAREA     1.4924 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.585 1.065 14.745 2.075 ;
        RECT  14.410 1.065 14.585 1.225 ;
        RECT  13.300 1.915 14.585 2.075 ;
        RECT  13.040 1.815 13.300 2.075 ;
        RECT  11.200 1.915 13.040 2.075 ;
        RECT  10.940 1.810 11.200 2.075 ;
        RECT  9.215 1.885 10.940 2.045 ;
        RECT  8.955 1.865 9.215 2.045 ;
        RECT  7.135 1.885 8.955 2.045 ;
        RECT  6.875 1.865 7.135 2.045 ;
        RECT  5.205 1.885 6.875 2.045 ;
        RECT  4.945 1.865 5.205 2.045 ;
        RECT  3.095 1.885 4.945 2.045 ;
        RECT  2.905 1.865 3.095 2.045 ;
        RECT  2.745 1.865 2.905 2.260 ;
        RECT  0.995 2.100 2.745 2.260 ;
        RECT  0.995 1.290 1.095 1.755 ;
        RECT  0.835 1.290 0.995 2.260 ;
        RECT  0.585 1.290 0.835 1.580 ;
        END
        ANTENNAGATEAREA     1.4924 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.145 1.460 14.405 1.705 ;
        RECT  13.630 1.460 14.145 1.620 ;
        RECT  13.560 1.385 13.630 1.620 ;
        RECT  13.350 1.385 13.560 1.630 ;
        RECT  10.680 1.470 13.350 1.630 ;
        RECT  10.470 1.470 10.680 1.705 ;
        RECT  10.420 1.525 10.470 1.705 ;
        RECT  9.890 1.525 10.420 1.685 ;
        RECT  9.630 1.525 9.890 1.705 ;
        RECT  6.675 1.525 9.630 1.685 ;
        RECT  6.390 1.525 6.675 1.705 ;
        RECT  2.515 1.525 6.390 1.685 ;
        RECT  2.355 1.525 2.515 1.920 ;
        RECT  1.695 1.760 2.355 1.920 ;
        RECT  1.695 1.290 1.715 1.580 ;
        RECT  1.535 1.290 1.695 1.920 ;
        RECT  1.505 1.290 1.535 1.730 ;
        RECT  1.315 1.470 1.505 1.730 ;
        END
        ANTENNAGATEAREA     1.4924 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.835 1.045 14.095 1.225 ;
        RECT  13.100 1.045 13.835 1.205 ;
        RECT  12.940 1.045 13.100 1.280 ;
        RECT  10.145 1.120 12.940 1.280 ;
        RECT  9.880 1.065 10.145 1.280 ;
        RECT  6.335 1.120 9.880 1.280 ;
        RECT  6.075 1.065 6.335 1.280 ;
        RECT  2.175 1.120 6.075 1.280 ;
        RECT  1.965 1.120 2.175 1.580 ;
        RECT  1.925 1.120 1.965 1.490 ;
        END
        ANTENNAGATEAREA     1.4924 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.395 -0.250 16.100 0.250 ;
        RECT  15.135 -0.250 15.395 0.405 ;
        RECT  14.300 -0.250 15.135 0.250 ;
        RECT  14.040 -0.250 14.300 0.405 ;
        RECT  13.220 -0.250 14.040 0.250 ;
        RECT  12.960 -0.250 13.220 0.405 ;
        RECT  12.140 -0.250 12.960 0.250 ;
        RECT  11.880 -0.250 12.140 0.405 ;
        RECT  11.060 -0.250 11.880 0.250 ;
        RECT  10.800 -0.250 11.060 0.405 ;
        RECT  9.980 -0.250 10.800 0.250 ;
        RECT  9.720 -0.250 9.980 0.405 ;
        RECT  8.895 -0.250 9.720 0.250 ;
        RECT  8.635 -0.250 8.895 0.405 ;
        RECT  7.815 -0.250 8.635 0.250 ;
        RECT  7.555 -0.250 7.815 0.405 ;
        RECT  6.735 -0.250 7.555 0.250 ;
        RECT  6.475 -0.250 6.735 0.405 ;
        RECT  5.655 -0.250 6.475 0.250 ;
        RECT  5.395 -0.250 5.655 0.405 ;
        RECT  4.575 -0.250 5.395 0.250 ;
        RECT  4.315 -0.250 4.575 0.405 ;
        RECT  3.495 -0.250 4.315 0.250 ;
        RECT  3.235 -0.250 3.495 0.405 ;
        RECT  2.415 -0.250 3.235 0.250 ;
        RECT  2.155 -0.250 2.415 0.405 ;
        RECT  1.325 -0.250 2.155 0.250 ;
        RECT  1.065 -0.250 1.325 0.405 ;
        RECT  0.385 -0.250 1.065 0.250 ;
        RECT  0.125 -0.250 0.385 1.135 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.735 3.440 16.100 3.940 ;
        RECT  15.475 3.285 15.735 3.940 ;
        RECT  11.905 3.440 15.475 3.940 ;
        RECT  11.645 3.285 11.905 3.940 ;
        RECT  7.820 3.440 11.645 3.940 ;
        RECT  7.560 3.285 7.820 3.940 ;
        RECT  3.800 3.440 7.560 3.940 ;
        RECT  3.540 3.285 3.800 3.940 ;
        RECT  0.585 3.440 3.540 3.940 ;
        RECT  0.325 2.945 0.585 3.940 ;
        RECT  0.000 3.440 0.325 3.940 ;
        END
    END VDD
END NOR4X8

MACRO NOR4X6
    CLASS CORE ;
    FOREIGN NOR4X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.960 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.640 0.470 11.835 3.105 ;
        RECT  11.625 0.470 11.640 1.355 ;
        RECT  11.625 2.745 11.640 3.105 ;
        RECT  11.165 0.470 11.625 1.170 ;
        RECT  1.835 2.815 11.625 3.105 ;
        RECT  10.695 0.880 11.165 1.170 ;
        RECT  10.340 0.585 10.695 1.170 ;
        RECT  0.955 0.585 10.340 0.875 ;
        RECT  0.665 0.585 0.955 1.110 ;
        END
        ANTENNADIFFAREA     3.0815 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.400 1.815 11.460 2.075 ;
        RECT  11.240 1.815 11.400 2.600 ;
        RECT  8.240 2.440 11.240 2.600 ;
        RECT  7.980 2.275 8.240 2.600 ;
        RECT  4.175 2.440 7.980 2.600 ;
        RECT  3.915 2.275 4.175 2.600 ;
        RECT  0.585 2.440 3.915 2.600 ;
        RECT  0.425 1.805 0.585 2.600 ;
        RECT  0.325 1.805 0.425 2.400 ;
        RECT  0.125 2.110 0.325 2.400 ;
        END
        ANTENNAGATEAREA     1.1050 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.060 1.385 11.200 1.545 ;
        RECT  10.900 1.385 11.060 2.095 ;
        RECT  9.215 1.935 10.900 2.095 ;
        RECT  8.955 1.815 9.215 2.095 ;
        RECT  7.135 1.935 8.955 2.095 ;
        RECT  6.875 1.815 7.135 2.095 ;
        RECT  5.205 1.935 6.875 2.095 ;
        RECT  4.945 1.810 5.205 2.095 ;
        RECT  3.095 1.935 4.945 2.095 ;
        RECT  2.995 1.810 3.095 2.095 ;
        RECT  2.835 1.810 2.995 2.260 ;
        RECT  1.095 2.100 2.835 2.260 ;
        RECT  0.935 1.290 1.095 2.260 ;
        RECT  0.835 1.290 0.935 1.755 ;
        RECT  0.585 1.290 0.835 1.580 ;
        END
        ANTENNAGATEAREA     1.1050 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.420 1.460 10.680 1.755 ;
        RECT  9.890 1.460 10.420 1.620 ;
        RECT  9.630 1.460 9.890 1.755 ;
        RECT  6.655 1.460 9.630 1.620 ;
        RECT  6.395 1.460 6.655 1.755 ;
        RECT  6.390 1.460 6.395 1.705 ;
        RECT  5.685 1.460 6.390 1.620 ;
        RECT  5.425 1.460 5.685 1.755 ;
        RECT  2.615 1.460 5.425 1.620 ;
        RECT  2.515 1.460 2.615 1.745 ;
        RECT  2.355 1.460 2.515 1.920 ;
        RECT  1.715 1.760 2.355 1.920 ;
        RECT  1.555 1.290 1.715 1.920 ;
        RECT  1.505 1.290 1.555 1.730 ;
        RECT  1.315 1.470 1.505 1.730 ;
        END
        ANTENNAGATEAREA     1.1050 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.880 1.065 10.145 1.280 ;
        RECT  6.335 1.120 9.880 1.280 ;
        RECT  6.075 1.065 6.335 1.280 ;
        RECT  2.175 1.120 6.075 1.280 ;
        RECT  1.965 1.120 2.175 1.580 ;
        RECT  1.925 1.120 1.965 1.385 ;
        END
        ANTENNAGATEAREA     1.1050 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.965 -0.250 11.960 0.250 ;
        RECT  10.705 -0.250 10.965 0.405 ;
        RECT  9.980 -0.250 10.705 0.250 ;
        RECT  9.720 -0.250 9.980 0.405 ;
        RECT  8.895 -0.250 9.720 0.250 ;
        RECT  8.635 -0.250 8.895 0.405 ;
        RECT  7.815 -0.250 8.635 0.250 ;
        RECT  7.555 -0.250 7.815 0.405 ;
        RECT  6.735 -0.250 7.555 0.250 ;
        RECT  6.475 -0.250 6.735 0.405 ;
        RECT  5.655 -0.250 6.475 0.250 ;
        RECT  5.395 -0.250 5.655 0.405 ;
        RECT  4.575 -0.250 5.395 0.250 ;
        RECT  4.315 -0.250 4.575 0.405 ;
        RECT  3.495 -0.250 4.315 0.250 ;
        RECT  3.235 -0.250 3.495 0.405 ;
        RECT  2.415 -0.250 3.235 0.250 ;
        RECT  2.155 -0.250 2.415 0.405 ;
        RECT  1.325 -0.250 2.155 0.250 ;
        RECT  1.065 -0.250 1.325 0.405 ;
        RECT  0.385 -0.250 1.065 0.250 ;
        RECT  0.125 -0.250 0.385 1.135 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.710 3.440 11.960 3.940 ;
        RECT  11.450 3.285 11.710 3.940 ;
        RECT  7.820 3.440 11.450 3.940 ;
        RECT  7.560 3.285 7.820 3.940 ;
        RECT  3.800 3.440 7.560 3.940 ;
        RECT  3.540 3.285 3.800 3.940 ;
        RECT  0.585 3.440 3.540 3.940 ;
        RECT  0.325 2.945 0.585 3.940 ;
        RECT  0.000 3.440 0.325 3.940 ;
        END
    END VDD
END NOR4X6

MACRO NOR4X4
    CLASS CORE ;
    FOREIGN NOR4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.530 0.585 7.710 3.105 ;
        RECT  7.485 0.585 7.530 1.580 ;
        RECT  5.915 2.875 7.530 3.105 ;
        RECT  6.195 0.585 7.485 0.785 ;
        RECT  5.935 0.495 6.195 0.785 ;
        RECT  5.115 0.585 5.935 0.785 ;
        RECT  5.655 2.875 5.915 3.155 ;
        RECT  2.065 2.875 5.655 3.105 ;
        RECT  4.855 0.495 5.115 0.785 ;
        RECT  4.035 0.585 4.855 0.785 ;
        RECT  3.775 0.495 4.035 0.785 ;
        RECT  2.955 0.585 3.775 0.785 ;
        RECT  2.695 0.495 2.955 0.785 ;
        RECT  1.875 0.585 2.695 0.785 ;
        RECT  1.805 2.875 2.065 3.135 ;
        RECT  1.615 0.495 1.875 0.785 ;
        RECT  0.925 0.585 1.615 0.785 ;
        RECT  0.765 0.585 0.925 1.110 ;
        RECT  0.665 0.850 0.765 1.110 ;
        END
        ANTENNADIFFAREA     2.0323 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.190 1.805 7.350 2.690 ;
        RECT  4.005 2.530 7.190 2.690 ;
        RECT  3.745 2.490 4.005 2.690 ;
        RECT  0.585 2.530 3.745 2.690 ;
        RECT  0.425 1.805 0.585 2.690 ;
        RECT  0.325 1.805 0.425 2.400 ;
        RECT  0.125 2.110 0.325 2.400 ;
        END
        ANTENNAGATEAREA     0.7293 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.960 1.325 7.090 1.585 ;
        RECT  6.800 1.325 6.960 2.310 ;
        RECT  4.940 2.150 6.800 2.310 ;
        RECT  4.655 1.645 4.940 2.310 ;
        RECT  3.095 2.150 4.655 2.310 ;
        RECT  2.835 1.810 3.095 2.310 ;
        RECT  0.995 2.150 2.835 2.310 ;
        RECT  0.995 1.290 1.095 1.755 ;
        RECT  0.835 1.290 0.995 2.310 ;
        RECT  0.585 1.290 0.835 1.580 ;
        END
        ANTENNAGATEAREA     0.7293 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.820 1.715 6.610 1.875 ;
        RECT  5.720 1.495 5.820 1.875 ;
        RECT  5.560 1.305 5.720 1.875 ;
        RECT  2.565 1.305 5.560 1.465 ;
        RECT  2.405 1.305 2.565 1.970 ;
        RECT  1.715 1.810 2.405 1.970 ;
        RECT  1.555 1.290 1.715 1.970 ;
        RECT  1.505 1.290 1.555 1.730 ;
        RECT  1.315 1.470 1.505 1.730 ;
        END
        ANTENNAGATEAREA     0.7293 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 1.185 6.535 1.445 ;
        RECT  6.275 0.965 6.435 1.445 ;
        RECT  2.175 0.965 6.275 1.125 ;
        RECT  2.085 0.965 2.175 1.580 ;
        RECT  2.015 0.965 2.085 1.630 ;
        RECT  1.965 1.290 2.015 1.630 ;
        RECT  1.925 1.370 1.965 1.630 ;
        END
        ANTENNAGATEAREA     0.7293 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.735 -0.250 7.820 0.250 ;
        RECT  6.475 -0.250 6.735 0.405 ;
        RECT  5.655 -0.250 6.475 0.250 ;
        RECT  5.395 -0.250 5.655 0.405 ;
        RECT  4.575 -0.250 5.395 0.250 ;
        RECT  4.315 -0.250 4.575 0.405 ;
        RECT  3.495 -0.250 4.315 0.250 ;
        RECT  3.235 -0.250 3.495 0.405 ;
        RECT  2.415 -0.250 3.235 0.250 ;
        RECT  2.155 -0.250 2.415 0.405 ;
        RECT  1.325 -0.250 2.155 0.250 ;
        RECT  1.065 -0.250 1.325 0.405 ;
        RECT  0.385 -0.250 1.065 0.250 ;
        RECT  0.125 -0.250 0.385 1.135 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.680 3.440 7.820 3.940 ;
        RECT  7.420 3.285 7.680 3.940 ;
        RECT  3.800 3.440 7.420 3.940 ;
        RECT  3.540 3.285 3.800 3.940 ;
        RECT  0.585 3.440 3.540 3.940 ;
        RECT  0.325 2.945 0.585 3.940 ;
        RECT  0.000 3.440 0.325 3.940 ;
        END
    END VDD
END NOR4X4

MACRO NOR4X2
    CLASS CORE ;
    FOREIGN NOR4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.355 0.850 3.615 1.110 ;
        RECT  2.705 0.900 3.355 1.060 ;
        RECT  2.445 0.430 2.705 1.060 ;
        RECT  2.425 0.695 2.445 1.060 ;
        RECT  1.785 0.900 2.425 1.060 ;
        RECT  0.265 2.820 2.205 2.980 ;
        RECT  1.715 0.800 1.785 1.060 ;
        RECT  1.685 0.695 1.715 1.060 ;
        RECT  1.525 0.585 1.685 1.060 ;
        RECT  0.785 0.585 1.525 0.745 ;
        RECT  0.625 0.585 0.785 1.115 ;
        RECT  0.585 0.695 0.625 1.115 ;
        RECT  0.335 0.855 0.585 1.115 ;
        RECT  0.265 0.855 0.335 1.170 ;
        RECT  0.105 0.855 0.265 2.980 ;
        END
        ANTENNADIFFAREA     1.3476 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.290 4.015 2.370 ;
        RECT  3.735 1.455 3.805 2.370 ;
        RECT  3.435 2.210 3.735 2.370 ;
        RECT  3.275 2.210 3.435 2.640 ;
        RECT  0.605 2.480 3.275 2.640 ;
        RECT  0.445 1.580 0.605 2.640 ;
        END
        ANTENNAGATEAREA     0.3848 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.475 1.515 3.555 1.990 ;
        RECT  3.215 1.290 3.475 2.030 ;
        RECT  3.045 1.870 3.215 2.030 ;
        RECT  2.885 1.870 3.045 2.300 ;
        RECT  1.255 2.140 2.885 2.300 ;
        RECT  1.135 1.925 1.255 2.300 ;
        RECT  0.975 1.270 1.135 2.300 ;
        RECT  0.925 1.270 0.975 1.530 ;
        END
        ANTENNAGATEAREA     0.3848 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.705 1.410 2.965 1.670 ;
        RECT  2.700 1.510 2.705 1.670 ;
        RECT  2.540 1.510 2.700 1.960 ;
        RECT  1.715 1.800 2.540 1.960 ;
        RECT  1.555 1.240 1.715 1.960 ;
        RECT  1.410 1.240 1.555 1.580 ;
        END
        ANTENNAGATEAREA     0.3848 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.240 2.355 1.620 ;
        END
        ANTENNAGATEAREA     0.3848 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 -0.250 4.140 0.250 ;
        RECT  3.755 -0.250 4.015 0.405 ;
        RECT  3.215 -0.250 3.755 0.250 ;
        RECT  2.955 -0.250 3.215 0.405 ;
        RECT  2.185 -0.250 2.955 0.250 ;
        RECT  1.925 -0.250 2.185 0.405 ;
        RECT  1.235 -0.250 1.925 0.250 ;
        RECT  0.975 -0.250 1.235 0.405 ;
        RECT  0.385 -0.250 0.975 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.550 4.015 3.940 ;
        RECT  0.385 3.440 3.755 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR4X2

MACRO NOR4X1
    CLASS CORE ;
    FOREIGN NOR4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.180 1.010 2.210 1.955 ;
        RECT  2.175 1.010 2.180 2.415 ;
        RECT  2.050 0.845 2.175 2.415 ;
        RECT  1.965 0.845 2.050 1.170 ;
        RECT  1.960 1.795 2.050 2.415 ;
        RECT  0.525 0.845 1.965 1.105 ;
        RECT  1.920 2.210 1.960 2.415 ;
        RECT  1.660 2.210 1.920 3.150 ;
        END
        ANTENNADIFFAREA     0.7417 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.525 0.370 1.985 ;
        RECT  0.125 1.525 0.335 1.990 ;
        RECT  0.090 1.525 0.125 1.985 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.290 0.875 1.550 ;
        RECT  0.585 1.290 0.835 1.820 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.340 1.440 1.500 ;
        RECT  1.230 1.700 1.255 1.990 ;
        RECT  1.065 1.340 1.230 1.990 ;
        RECT  1.045 1.700 1.065 1.990 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.780 1.350 1.870 1.610 ;
        RECT  1.715 1.350 1.780 1.930 ;
        RECT  1.620 1.350 1.715 1.990 ;
        RECT  1.505 1.700 1.620 1.990 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.135 -0.250 2.300 0.250 ;
        RECT  1.875 -0.250 2.135 0.405 ;
        RECT  1.185 -0.250 1.875 0.250 ;
        RECT  0.925 -0.250 1.185 0.405 ;
        RECT  0.385 -0.250 0.925 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.450 3.440 2.300 3.940 ;
        RECT  0.190 2.215 0.450 3.940 ;
        RECT  0.000 3.440 0.190 3.940 ;
        END
    END VDD
END NOR4X1

MACRO NOR4XL
    CLASS CORE ;
    FOREIGN NOR4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.690 2.180 2.040 2.440 ;
        RECT  1.675 0.915 1.935 1.085 ;
        RECT  0.795 2.180 1.690 2.340 ;
        RECT  0.685 0.925 1.675 1.085 ;
        RECT  0.685 2.110 0.795 2.400 ;
        RECT  0.585 0.925 0.685 2.400 ;
        RECT  0.525 0.925 0.585 2.335 ;
        RECT  0.410 0.990 0.525 1.250 ;
        END
        ANTENNADIFFAREA     0.6553 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.330 1.700 0.335 1.990 ;
        RECT  0.090 1.645 0.330 2.165 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 1.515 1.255 1.990 ;
        RECT  1.045 1.360 1.160 1.990 ;
        RECT  1.000 1.360 1.045 1.925 ;
        RECT  0.865 1.360 1.000 1.635 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.510 1.265 1.725 1.735 ;
        RECT  1.435 1.265 1.510 1.635 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.165 1.515 2.175 1.990 ;
        RECT  1.955 1.320 2.165 1.990 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 -0.250 2.300 0.250 ;
        RECT  1.675 -0.250 1.935 0.405 ;
        RECT  1.360 -0.250 1.675 0.250 ;
        RECT  1.100 -0.250 1.360 0.405 ;
        RECT  0.580 -0.250 1.100 0.250 ;
        RECT  0.320 -0.250 0.580 0.405 ;
        RECT  0.000 -0.250 0.320 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.565 3.440 2.300 3.940 ;
        RECT  0.305 2.605 0.565 3.940 ;
        RECT  0.000 3.440 0.305 3.940 ;
        END
    END VDD
END NOR4XL

MACRO NOR3X8
    CLASS CORE ;
    FOREIGN NOR3X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.595 0.585 9.075 2.995 ;
        RECT  1.205 0.585 8.595 0.800 ;
        RECT  8.405 2.110 8.595 2.995 ;
        RECT  6.330 2.595 8.405 2.995 ;
        RECT  6.070 2.595 6.330 3.195 ;
        RECT  4.005 2.595 6.070 2.995 ;
        RECT  3.745 2.595 4.005 3.195 ;
        RECT  1.685 2.595 3.745 2.995 ;
        RECT  1.425 2.595 1.685 3.195 ;
        RECT  0.945 0.585 1.205 0.910 ;
        END
        ANTENNADIFFAREA     3.1859 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.320 1.660 7.465 1.820 ;
        RECT  7.160 1.660 7.320 2.330 ;
        RECT  5.395 2.170 7.160 2.330 ;
        RECT  5.370 1.925 5.395 2.330 ;
        RECT  5.110 1.665 5.370 2.330 ;
        RECT  4.910 2.110 5.110 2.330 ;
        RECT  2.645 2.170 4.910 2.330 ;
        RECT  2.380 1.665 2.645 2.330 ;
        RECT  0.610 2.170 2.380 2.330 ;
        RECT  0.555 2.110 0.610 2.330 ;
        RECT  0.395 1.575 0.555 2.330 ;
        RECT  0.295 1.575 0.395 1.990 ;
        RECT  0.125 1.700 0.295 1.990 ;
        END
        ANTENNAGATEAREA     1.3520 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.850 1.405 7.945 1.665 ;
        RECT  7.685 1.320 7.850 1.665 ;
        RECT  6.980 1.320 7.685 1.480 ;
        RECT  6.820 1.320 6.980 1.920 ;
        RECT  6.720 1.615 6.820 1.920 ;
        RECT  5.850 1.760 6.720 1.920 ;
        RECT  5.690 1.325 5.850 1.920 ;
        RECT  5.590 1.325 5.690 1.490 ;
        RECT  4.750 1.325 5.590 1.485 ;
        RECT  4.545 1.325 4.750 1.490 ;
        RECT  4.385 1.325 4.545 1.750 ;
        RECT  3.215 1.590 4.385 1.750 ;
        RECT  3.055 1.325 3.215 1.750 ;
        RECT  2.955 1.325 3.055 1.505 ;
        RECT  2.175 1.325 2.955 1.485 ;
        RECT  1.965 1.325 2.175 1.990 ;
        RECT  1.905 1.325 1.965 1.880 ;
        RECT  1.035 1.720 1.905 1.880 ;
        RECT  0.775 1.595 1.035 1.880 ;
        END
        ANTENNAGATEAREA     1.3520 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.215 0.980 8.375 1.585 ;
        RECT  6.330 0.980 8.215 1.140 ;
        RECT  6.105 0.980 6.330 1.580 ;
        RECT  6.070 0.980 6.105 1.515 ;
        RECT  4.175 0.980 6.070 1.140 ;
        RECT  3.575 0.980 4.175 1.405 ;
        RECT  1.545 0.980 3.575 1.140 ;
        RECT  1.385 0.980 1.545 1.535 ;
        RECT  1.285 1.275 1.385 1.535 ;
        END
        ANTENNAGATEAREA     1.3520 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.265 -0.250 9.200 0.250 ;
        RECT  8.005 -0.250 8.265 0.405 ;
        RECT  7.185 -0.250 8.005 0.250 ;
        RECT  6.925 -0.250 7.185 0.405 ;
        RECT  6.100 -0.250 6.925 0.250 ;
        RECT  5.840 -0.250 6.100 0.405 ;
        RECT  5.015 -0.250 5.840 0.250 ;
        RECT  4.755 -0.250 5.015 0.405 ;
        RECT  3.925 -0.250 4.755 0.250 ;
        RECT  3.665 -0.250 3.925 0.405 ;
        RECT  2.845 -0.250 3.665 0.250 ;
        RECT  2.585 -0.250 2.845 0.405 ;
        RECT  1.750 -0.250 2.585 0.250 ;
        RECT  1.490 -0.250 1.750 0.405 ;
        RECT  0.660 -0.250 1.490 0.250 ;
        RECT  0.400 -0.250 0.660 1.145 ;
        RECT  0.000 -0.250 0.400 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.665 3.440 9.200 3.940 ;
        RECT  7.405 3.285 7.665 3.940 ;
        RECT  5.170 3.440 7.405 3.940 ;
        RECT  4.910 3.285 5.170 3.940 ;
        RECT  2.845 3.440 4.910 3.940 ;
        RECT  2.585 3.285 2.845 3.940 ;
        RECT  0.385 3.440 2.585 3.940 ;
        RECT  0.125 2.590 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR3X8

MACRO NOR3X6
    CLASS CORE ;
    FOREIGN NOR3X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.940 0.590 7.240 3.220 ;
        RECT  6.645 0.590 6.940 0.890 ;
        RECT  6.565 2.520 6.940 3.220 ;
        RECT  6.385 0.590 6.645 1.090 ;
        RECT  6.330 2.595 6.565 2.895 ;
        RECT  1.205 0.590 6.385 0.775 ;
        RECT  6.070 2.595 6.330 3.195 ;
        RECT  4.015 2.595 6.070 2.895 ;
        RECT  4.005 2.595 4.015 2.995 ;
        RECT  3.745 2.595 4.005 3.195 ;
        RECT  3.530 2.595 3.745 3.045 ;
        RECT  1.405 2.745 3.530 3.045 ;
        RECT  0.945 0.590 1.205 0.910 ;
        END
        ANTENNADIFFAREA     2.6907 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.600 1.600 6.760 2.250 ;
        RECT  5.395 2.090 6.600 2.250 ;
        RECT  5.370 1.925 5.395 2.250 ;
        RECT  5.105 1.635 5.370 2.250 ;
        RECT  2.645 2.090 5.105 2.250 ;
        RECT  2.540 1.635 2.645 2.250 ;
        RECT  2.380 1.635 2.540 2.505 ;
        RECT  0.555 2.345 2.380 2.505 ;
        RECT  0.395 1.575 0.555 2.505 ;
        RECT  0.295 1.575 0.395 1.990 ;
        RECT  0.125 1.700 0.295 1.990 ;
        END
        ANTENNAGATEAREA     1.1180 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.590 1.295 5.850 1.475 ;
        RECT  4.645 1.295 5.590 1.455 ;
        RECT  4.545 1.295 4.645 1.470 ;
        RECT  4.385 1.295 4.545 1.910 ;
        RECT  3.215 1.750 4.385 1.910 ;
        RECT  3.055 1.295 3.215 1.910 ;
        RECT  2.125 1.295 3.055 1.455 ;
        RECT  2.125 1.700 2.175 1.990 ;
        RECT  1.965 1.295 2.125 2.165 ;
        RECT  1.765 1.295 1.965 1.455 ;
        RECT  1.035 2.005 1.965 2.165 ;
        RECT  0.875 1.580 1.035 2.165 ;
        RECT  0.775 1.580 0.875 1.840 ;
        END
        ANTENNAGATEAREA     1.1180 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 1.405 6.330 1.665 ;
        RECT  6.190 1.290 6.315 1.665 ;
        RECT  6.070 0.955 6.190 1.665 ;
        RECT  6.030 0.955 6.070 1.615 ;
        RECT  3.955 0.955 6.030 1.115 ;
        RECT  3.695 0.955 3.955 1.395 ;
        RECT  1.545 0.955 3.695 1.115 ;
        RECT  1.385 0.955 1.545 1.825 ;
        RECT  1.285 1.565 1.385 1.825 ;
        END
        ANTENNAGATEAREA     1.1180 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 -0.250 7.360 0.250 ;
        RECT  6.925 -0.250 7.185 0.405 ;
        RECT  6.100 -0.250 6.925 0.250 ;
        RECT  5.840 -0.250 6.100 0.405 ;
        RECT  5.015 -0.250 5.840 0.250 ;
        RECT  4.755 -0.250 5.015 0.405 ;
        RECT  3.925 -0.250 4.755 0.250 ;
        RECT  3.665 -0.250 3.925 0.405 ;
        RECT  2.845 -0.250 3.665 0.250 ;
        RECT  2.585 -0.250 2.845 0.405 ;
        RECT  1.750 -0.250 2.585 0.250 ;
        RECT  1.490 -0.250 1.750 0.405 ;
        RECT  0.665 -0.250 1.490 0.250 ;
        RECT  0.405 -0.250 0.665 1.145 ;
        RECT  0.000 -0.250 0.405 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.170 3.440 7.360 3.940 ;
        RECT  4.910 3.285 5.170 3.940 ;
        RECT  2.845 3.440 4.910 3.940 ;
        RECT  2.585 3.285 2.845 3.940 ;
        RECT  0.385 3.440 2.585 3.940 ;
        RECT  0.125 2.865 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR3X6

MACRO NOR3X4
    CLASS CORE ;
    FOREIGN NOR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.390 1.105 5.395 2.810 ;
        RECT  5.385 1.105 5.390 2.885 ;
        RECT  5.185 0.920 5.385 2.885 ;
        RECT  3.830 0.920 5.185 1.120 ;
        RECT  3.835 2.685 5.185 2.885 ;
        RECT  3.530 2.625 3.835 2.885 ;
        RECT  3.755 0.880 3.830 1.120 ;
        RECT  3.495 0.520 3.755 1.120 ;
        RECT  1.515 2.685 3.530 2.885 ;
        RECT  1.595 0.605 3.495 0.805 ;
        RECT  1.335 0.575 1.595 0.835 ;
        RECT  1.255 2.625 1.515 2.885 ;
        END
        ANTENNADIFFAREA     1.6560 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 1.700 4.935 2.175 ;
        RECT  4.785 1.680 4.885 2.175 ;
        RECT  4.625 1.680 4.785 2.360 ;
        RECT  4.450 2.110 4.625 2.360 ;
        RECT  2.545 2.200 4.450 2.360 ;
        RECT  2.385 1.670 2.545 2.360 ;
        RECT  0.795 2.200 2.385 2.360 ;
        RECT  0.755 1.925 0.795 2.360 ;
        RECT  0.585 1.645 0.755 2.360 ;
        RECT  0.295 1.645 0.585 1.805 ;
        END
        ANTENNAGATEAREA     0.7540 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.145 1.305 4.405 1.565 ;
        RECT  3.225 1.355 4.145 1.515 ;
        RECT  3.065 0.985 3.225 1.515 ;
        RECT  1.865 0.985 3.065 1.145 ;
        RECT  1.705 0.985 1.865 1.545 ;
        RECT  1.605 1.280 1.705 1.545 ;
        RECT  0.590 1.280 1.605 1.440 ;
        RECT  0.335 1.115 0.590 1.440 ;
        RECT  0.170 0.880 0.335 1.440 ;
        RECT  0.125 0.880 0.170 1.170 ;
        END
        ANTENNAGATEAREA     0.7540 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.700 4.015 1.990 ;
        RECT  3.530 1.715 3.805 1.990 ;
        RECT  2.910 1.830 3.530 1.990 ;
        RECT  2.885 1.765 2.910 1.990 ;
        RECT  2.725 1.330 2.885 1.990 ;
        RECT  2.205 1.330 2.725 1.490 ;
        RECT  2.045 1.330 2.205 2.015 ;
        RECT  1.345 1.855 2.045 2.015 ;
        RECT  1.185 1.645 1.345 2.015 ;
        RECT  1.085 1.645 1.185 1.805 ;
        END
        ANTENNAGATEAREA     0.7540 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.295 -0.250 5.520 0.250 ;
        RECT  4.035 -0.250 4.295 0.405 ;
        RECT  3.215 -0.250 4.035 0.250 ;
        RECT  2.955 -0.250 3.215 0.405 ;
        RECT  2.135 -0.250 2.955 0.250 ;
        RECT  1.875 -0.250 2.135 0.405 ;
        RECT  1.045 -0.250 1.875 0.250 ;
        RECT  0.785 -0.250 1.045 1.095 ;
        RECT  0.000 -0.250 0.785 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.060 3.440 5.520 3.940 ;
        RECT  4.800 3.285 5.060 3.940 ;
        RECT  2.675 3.440 4.800 3.940 ;
        RECT  2.415 3.285 2.675 3.940 ;
        RECT  0.385 3.440 2.415 3.940 ;
        RECT  0.125 2.075 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR3X4

MACRO NOR3X2
    CLASS CORE ;
    FOREIGN NOR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 0.695 2.635 0.945 ;
        RECT  2.425 0.585 2.585 1.435 ;
        RECT  1.990 0.585 2.425 0.745 ;
        RECT  2.055 1.275 2.425 1.435 ;
        RECT  1.895 1.275 2.055 2.330 ;
        RECT  1.725 0.545 1.990 0.745 ;
        RECT  1.520 2.170 1.895 2.330 ;
        RECT  0.900 0.585 1.725 0.745 ;
        RECT  1.260 2.170 1.520 2.430 ;
        RECT  0.795 0.495 0.900 1.095 ;
        RECT  0.640 0.470 0.795 1.095 ;
        RECT  0.585 0.470 0.640 0.945 ;
        END
        ANTENNADIFFAREA     0.8359 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.495 1.700 2.635 1.990 ;
        RECT  2.395 1.620 2.495 1.990 ;
        RECT  2.235 1.620 2.395 2.770 ;
        RECT  2.150 2.520 2.235 2.770 ;
        RECT  0.795 2.610 2.150 2.770 ;
        RECT  0.730 1.925 0.795 2.770 ;
        RECT  0.570 1.500 0.730 2.770 ;
        RECT  0.560 1.500 0.570 1.660 ;
        RECT  0.300 1.400 0.560 1.660 ;
        END
        ANTENNAGATEAREA     0.3458 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 0.935 2.245 1.095 ;
        RECT  1.555 0.935 1.715 1.390 ;
        RECT  1.255 1.230 1.555 1.390 ;
        RECT  1.080 1.230 1.255 1.580 ;
        RECT  1.045 1.290 1.080 1.580 ;
        RECT  0.960 1.315 1.045 1.550 ;
        RECT  0.910 1.315 0.960 1.475 ;
        END
        ANTENNAGATEAREA     0.3458 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 1.700 1.715 1.990 ;
        RECT  1.480 1.570 1.640 1.990 ;
        RECT  1.295 1.760 1.480 1.990 ;
        END
        ANTENNAGATEAREA     0.3458 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 -0.250 2.760 0.250 ;
        RECT  1.185 -0.250 1.445 0.405 ;
        RECT  0.390 -0.250 1.185 0.250 ;
        RECT  0.130 -0.250 0.390 1.110 ;
        RECT  0.000 -0.250 0.130 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 3.440 2.760 3.940 ;
        RECT  2.375 3.285 2.635 3.940 ;
        RECT  0.390 3.440 2.375 3.940 ;
        RECT  0.130 1.955 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
END NOR3X2

MACRO NOR3X1
    CLASS CORE ;
    FOREIGN NOR3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 0.435 1.715 1.105 ;
        RECT  1.545 2.745 1.715 2.995 ;
        RECT  1.285 2.255 1.545 3.195 ;
        RECT  1.445 0.435 1.505 0.595 ;
        RECT  0.700 0.945 1.505 1.105 ;
        RECT  0.795 2.255 1.285 2.415 ;
        RECT  0.700 2.110 0.795 2.415 ;
        RECT  0.660 0.945 0.700 2.415 ;
        RECT  0.585 0.845 0.660 2.415 ;
        RECT  0.540 0.845 0.585 2.360 ;
        RECT  0.400 0.845 0.540 1.105 ;
        END
        ANTENNADIFFAREA     0.8724 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.320 1.290 0.335 1.765 ;
        RECT  0.160 1.290 0.320 2.135 ;
        RECT  0.125 1.290 0.160 1.765 ;
        END
        ANTENNAGATEAREA     0.1755 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.035 1.290 1.280 1.825 ;
        RECT  0.880 1.565 1.035 1.825 ;
        END
        ANTENNAGATEAREA     0.1755 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.510 1.715 2.000 ;
        END
        ANTENNAGATEAREA     0.1755 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 -0.250 1.840 0.250 ;
        RECT  0.590 -0.250 1.190 0.405 ;
        RECT  0.000 -0.250 0.590 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 1.840 3.940 ;
        RECT  0.125 2.540 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR3X1

MACRO NOR3XL
    CLASS CORE ;
    FOREIGN NOR3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.535 0.880 1.715 2.425 ;
        RECT  1.530 0.880 1.535 1.355 ;
        RECT  1.435 2.165 1.535 2.425 ;
        RECT  1.505 0.880 1.530 1.295 ;
        RECT  1.395 1.035 1.505 1.295 ;
        RECT  0.645 1.065 1.395 1.225 ;
        RECT  0.385 1.015 0.645 1.275 ;
        END
        ANTENNADIFFAREA     0.5358 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.545 0.395 2.030 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 1.455 0.925 1.615 ;
        RECT  0.795 1.455 0.840 1.935 ;
        RECT  0.585 1.455 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.725 1.355 1.985 ;
        RECT  1.095 1.725 1.255 2.400 ;
        RECT  1.045 2.110 1.095 2.400 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.225 -0.250 1.840 0.250 ;
        RECT  0.965 -0.250 1.225 0.795 ;
        RECT  0.645 -0.250 0.965 0.250 ;
        RECT  0.385 -0.250 0.645 0.405 ;
        RECT  0.000 -0.250 0.385 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 1.840 3.940 ;
        RECT  0.125 2.215 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR3XL

MACRO NOR2X8
    CLASS CORE ;
    FOREIGN NOR2X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.905 0.585 5.395 2.810 ;
        RECT  4.585 0.585 4.905 1.095 ;
        RECT  4.725 2.110 4.905 2.810 ;
        RECT  4.485 2.275 4.725 2.810 ;
        RECT  4.325 0.495 4.585 1.095 ;
        RECT  4.225 2.275 4.485 3.215 ;
        RECT  3.505 0.585 4.325 0.985 ;
        RECT  2.910 2.275 4.225 2.675 ;
        RECT  3.245 0.495 3.505 1.095 ;
        RECT  2.425 0.585 3.245 0.985 ;
        RECT  2.845 2.275 2.910 2.810 ;
        RECT  2.585 2.275 2.845 3.215 ;
        RECT  2.425 2.275 2.585 2.995 ;
        RECT  2.165 0.495 2.425 1.095 ;
        RECT  1.255 2.275 2.425 2.675 ;
        RECT  1.345 0.585 2.165 0.985 ;
        RECT  1.085 0.495 1.345 1.095 ;
        RECT  1.205 2.275 1.255 2.995 ;
        RECT  0.945 2.275 1.205 3.215 ;
        END
        ANTENNADIFFAREA     2.6764 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.545 1.635 3.645 1.795 ;
        RECT  3.385 1.635 3.545 1.985 ;
        RECT  2.195 1.825 3.385 1.985 ;
        RECT  1.595 1.630 2.195 1.985 ;
        RECT  0.555 1.825 1.595 1.985 ;
        RECT  0.335 1.585 0.555 1.985 ;
        RECT  0.295 1.585 0.335 1.990 ;
        RECT  0.125 1.700 0.295 1.990 ;
        END
        ANTENNAGATEAREA     1.2714 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.560 4.725 1.820 ;
        RECT  4.450 1.560 4.475 1.990 ;
        RECT  4.425 1.515 4.450 1.990 ;
        RECT  4.265 1.275 4.425 1.990 ;
        RECT  3.015 1.275 4.265 1.455 ;
        RECT  2.415 1.275 3.015 1.645 ;
        RECT  1.145 1.275 2.415 1.435 ;
        RECT  0.985 1.275 1.145 1.645 ;
        RECT  0.775 1.385 0.985 1.645 ;
        END
        ANTENNAGATEAREA     1.2714 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.125 -0.250 5.520 0.250 ;
        RECT  4.865 -0.250 5.125 0.405 ;
        RECT  4.045 -0.250 4.865 0.250 ;
        RECT  3.785 -0.250 4.045 0.405 ;
        RECT  2.965 -0.250 3.785 0.250 ;
        RECT  2.705 -0.250 2.965 0.405 ;
        RECT  1.885 -0.250 2.705 0.250 ;
        RECT  1.625 -0.250 1.885 0.405 ;
        RECT  0.805 -0.250 1.625 0.250 ;
        RECT  0.545 -0.250 0.805 1.145 ;
        RECT  0.000 -0.250 0.545 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.665 3.440 5.520 3.940 ;
        RECT  3.405 2.955 3.665 3.940 ;
        RECT  2.025 3.440 3.405 3.940 ;
        RECT  1.765 2.955 2.025 3.940 ;
        RECT  0.385 3.440 1.765 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR2X8

MACRO NOR2X6
    CLASS CORE ;
    FOREIGN NOR2X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.715 0.780 4.015 2.810 ;
        RECT  3.530 0.780 3.715 1.170 ;
        RECT  3.345 2.110 3.715 2.810 ;
        RECT  1.655 0.780 3.530 1.080 ;
        RECT  2.910 2.285 3.345 2.585 ;
        RECT  2.595 2.285 2.910 3.020 ;
        RECT  1.255 2.285 2.595 2.585 ;
        RECT  1.070 0.865 1.655 1.080 ;
        RECT  0.955 2.285 1.255 3.020 ;
        RECT  0.895 0.865 1.070 1.095 ;
        RECT  0.635 0.495 0.895 1.095 ;
        RECT  0.585 0.695 0.635 0.945 ;
        END
        ANTENNADIFFAREA     1.7856 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.265 1.385 3.525 1.645 ;
        RECT  3.095 1.485 3.265 1.645 ;
        RECT  2.935 1.485 3.095 2.025 ;
        RECT  2.225 1.865 2.935 2.025 ;
        RECT  1.965 1.600 2.225 2.025 ;
        RECT  0.795 1.865 1.965 2.025 ;
        RECT  0.770 1.700 0.795 2.025 ;
        RECT  0.610 1.655 0.770 2.025 ;
        RECT  0.585 1.655 0.610 1.990 ;
        RECT  0.520 1.655 0.585 1.815 ;
        RECT  0.260 1.555 0.520 1.815 ;
        END
        ANTENNAGATEAREA     0.9048 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.390 2.705 1.650 ;
        RECT  2.610 1.290 2.635 1.650 ;
        RECT  2.445 1.260 2.610 1.650 ;
        RECT  2.425 1.260 2.445 1.580 ;
        RECT  1.780 1.260 2.425 1.420 ;
        RECT  1.620 1.260 1.780 1.585 ;
        RECT  1.405 1.425 1.620 1.585 ;
        RECT  1.145 1.425 1.405 1.685 ;
        END
        ANTENNAGATEAREA     0.9048 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.535 -0.250 4.140 0.250 ;
        RECT  3.275 -0.250 3.535 0.405 ;
        RECT  2.455 -0.250 3.275 0.250 ;
        RECT  2.195 -0.250 2.455 0.405 ;
        RECT  1.405 -0.250 2.195 0.250 ;
        RECT  1.145 -0.250 1.405 0.685 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.190 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.725 3.440 4.140 3.940 ;
        RECT  3.465 3.285 3.725 3.940 ;
        RECT  2.055 3.440 3.465 3.940 ;
        RECT  1.795 2.790 2.055 3.940 ;
        RECT  0.385 3.440 1.795 3.940 ;
        RECT  0.125 2.215 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR2X6

MACRO NOR2X4
    CLASS CORE ;
    FOREIGN NOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 0.985 3.095 3.180 ;
        RECT  2.020 0.985 2.885 1.185 ;
        RECT  2.745 2.200 2.885 3.180 ;
        RECT  1.365 2.200 2.745 2.400 ;
        RECT  1.790 0.510 2.020 1.185 ;
        RECT  1.760 0.510 1.790 1.170 ;
        RECT  1.690 0.880 1.760 1.170 ;
        RECT  0.940 0.910 1.690 1.110 ;
        RECT  1.105 2.200 1.365 2.970 ;
        RECT  0.680 0.510 0.940 1.110 ;
        RECT  0.585 0.695 0.680 0.945 ;
        END
        ANTENNADIFFAREA     1.4703 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.755 1.730 2.015 1.990 ;
        RECT  0.610 1.795 1.755 1.955 ;
        RECT  0.595 1.765 0.610 1.955 ;
        RECT  0.335 1.405 0.595 1.955 ;
        RECT  0.125 1.700 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.6552 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.410 1.380 2.670 1.670 ;
        RECT  1.280 1.380 2.410 1.540 ;
        RECT  1.255 1.380 1.280 1.615 ;
        RECT  1.045 1.290 1.255 1.615 ;
        RECT  1.020 1.455 1.045 1.615 ;
        END
        ANTENNAGATEAREA     0.6552 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 -0.250 3.220 0.250 ;
        RECT  2.560 0.535 2.900 0.795 ;
        RECT  2.300 -0.250 2.560 0.795 ;
        RECT  1.480 -0.250 2.300 0.250 ;
        RECT  1.220 -0.250 1.480 0.405 ;
        RECT  0.385 -0.250 1.220 0.250 ;
        RECT  0.125 -0.250 0.385 1.170 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.185 3.440 3.220 3.940 ;
        RECT  1.925 2.580 2.185 3.940 ;
        RECT  0.495 3.440 1.925 3.940 ;
        RECT  0.235 2.210 0.495 3.940 ;
        RECT  0.000 3.440 0.235 3.940 ;
        END
    END VDD
END NOR2X4

MACRO NOR2X2
    CLASS CORE ;
    FOREIGN NOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 1.290 2.175 1.765 ;
        RECT  1.965 0.980 2.125 2.020 ;
        RECT  1.515 0.980 1.965 1.140 ;
        RECT  1.675 1.860 1.965 2.020 ;
        RECT  1.515 1.860 1.675 2.475 ;
        RECT  1.255 0.540 1.515 1.140 ;
        RECT  1.265 2.315 1.515 2.475 ;
        RECT  1.005 2.315 1.265 2.915 ;
        END
        ANTENNADIFFAREA     0.6384 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 1.360 1.745 1.680 ;
        RECT  0.485 1.360 1.485 1.520 ;
        RECT  0.325 1.360 0.485 2.005 ;
        RECT  0.225 1.700 0.325 2.005 ;
        RECT  0.125 1.700 0.225 1.990 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.150 1.700 1.255 1.990 ;
        RECT  1.045 1.700 1.150 2.095 ;
        RECT  0.850 1.705 1.045 2.095 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.055 -0.250 2.300 0.250 ;
        RECT  1.795 -0.250 2.055 0.800 ;
        RECT  0.975 -0.250 1.795 0.250 ;
        RECT  0.715 -0.250 0.975 1.140 ;
        RECT  0.000 -0.250 0.715 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 3.440 2.300 3.940 ;
        RECT  1.855 2.210 2.115 3.940 ;
        RECT  0.415 3.440 1.855 3.940 ;
        RECT  0.155 2.215 0.415 3.940 ;
        RECT  0.000 3.440 0.155 3.940 ;
        END
    END VDD
END NOR2X2

MACRO NOR2X1
    CLASS CORE ;
    FOREIGN NOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.380 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.095 0.880 1.255 2.775 ;
        RECT  1.045 0.880 1.095 1.170 ;
        RECT  0.905 2.175 1.095 2.775 ;
        RECT  0.825 0.880 1.045 1.095 ;
        RECT  0.565 0.835 0.825 1.095 ;
        END
        ANTENNADIFFAREA     0.4452 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.500 0.405 2.000 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.425 0.915 1.685 ;
        RECT  0.585 1.425 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 -0.250 1.380 0.250 ;
        RECT  0.245 -0.250 1.185 0.405 ;
        RECT  0.000 -0.250 0.245 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 1.380 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR2X1

MACRO NOR2XL
    CLASS CORE ;
    FOREIGN NOR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.380 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 2.110 1.255 2.400 ;
        RECT  1.070 1.135 1.230 2.460 ;
        RECT  0.815 1.135 1.070 1.295 ;
        RECT  1.045 2.110 1.070 2.460 ;
        RECT  0.835 2.200 1.045 2.460 ;
        RECT  0.555 1.035 0.815 1.295 ;
        END
        ANTENNADIFFAREA     0.2738 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.120 1.500 0.390 2.005 ;
        END
        ANTENNAGATEAREA     0.0871 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.565 0.875 1.990 ;
        END
        ANTENNAGATEAREA     0.0871 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 -0.250 1.380 0.250 ;
        RECT  0.985 -0.250 1.245 0.405 ;
        RECT  0.395 -0.250 0.985 0.250 ;
        RECT  0.135 -0.250 0.395 0.405 ;
        RECT  0.000 -0.250 0.135 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 1.380 3.940 ;
        RECT  0.125 2.890 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NOR2XL

MACRO NAND4BBX4
    CLASS CORE ;
    FOREIGN NAND4BBX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.595 0.695 8.615 3.080 ;
        RECT  8.355 0.615 8.595 3.080 ;
        RECT  5.705 0.615 8.355 0.855 ;
        RECT  1.295 2.820 8.355 3.080 ;
        RECT  5.445 0.505 5.705 1.105 ;
        RECT  3.800 0.865 5.445 1.105 ;
        RECT  3.530 0.855 3.800 1.105 ;
        RECT  2.760 0.855 3.530 1.095 ;
        RECT  2.500 0.495 2.760 1.095 ;
        END
        ANTENNADIFFAREA     2.5698 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.150 1.700 7.235 2.175 ;
        RECT  7.050 1.615 7.150 2.175 ;
        RECT  6.890 1.615 7.050 2.615 ;
        RECT  1.260 2.455 6.890 2.615 ;
        RECT  1.100 1.595 1.260 2.615 ;
        RECT  1.045 1.595 1.100 2.175 ;
        RECT  1.000 1.595 1.045 1.855 ;
        END
        ANTENNAGATEAREA     0.7098 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 1.615 6.665 1.875 ;
        RECT  6.405 1.615 6.565 2.275 ;
        RECT  4.740 2.115 6.405 2.275 ;
        RECT  4.480 2.025 4.740 2.275 ;
        RECT  3.780 2.025 4.480 2.185 ;
        RECT  3.520 2.025 3.780 2.275 ;
        RECT  1.740 2.115 3.520 2.275 ;
        RECT  1.580 1.615 1.740 2.275 ;
        RECT  1.505 1.615 1.580 1.990 ;
        RECT  1.480 1.615 1.505 1.875 ;
        END
        ANTENNAGATEAREA     0.7098 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.480 1.595 7.695 2.465 ;
        RECT  7.435 1.595 7.480 1.855 ;
        END
        ANTENNAGATEAREA     0.2743 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.730 1.925 0.795 2.400 ;
        RECT  0.570 1.595 0.730 2.400 ;
        END
        ANTENNAGATEAREA     0.2743 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.380 -0.250 8.740 0.250 ;
        RECT  7.120 -0.250 7.380 0.405 ;
        RECT  4.260 -0.250 7.120 0.250 ;
        RECT  4.000 -0.250 4.260 0.685 ;
        RECT  1.200 -0.250 4.000 0.250 ;
        RECT  0.940 -0.250 1.200 1.075 ;
        RECT  0.000 -0.250 0.940 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.500 3.440 8.740 3.940 ;
        RECT  7.240 3.285 7.500 3.940 ;
        RECT  6.415 3.440 7.240 3.940 ;
        RECT  6.155 3.285 6.415 3.940 ;
        RECT  5.330 3.440 6.155 3.940 ;
        RECT  4.730 3.285 5.330 3.940 ;
        RECT  3.530 3.440 4.730 3.940 ;
        RECT  2.930 3.285 3.530 3.940 ;
        RECT  2.110 3.440 2.930 3.940 ;
        RECT  1.850 3.285 2.110 3.940 ;
        RECT  1.020 3.440 1.850 3.940 ;
        RECT  0.760 2.935 1.020 3.940 ;
        RECT  0.000 3.440 0.760 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.035 1.965 8.135 2.565 ;
        RECT  7.875 1.065 8.035 2.565 ;
        RECT  6.190 1.065 7.875 1.225 ;
        RECT  6.030 1.065 6.190 1.935 ;
        RECT  5.925 1.615 6.030 1.935 ;
        RECT  5.220 1.775 5.925 1.935 ;
        RECT  5.440 1.285 5.700 1.545 ;
        RECT  2.820 1.285 5.440 1.445 ;
        RECT  4.960 1.665 5.220 1.935 ;
        RECT  3.320 1.665 4.960 1.825 ;
        RECT  3.040 1.665 3.320 1.895 ;
        RECT  2.220 1.735 3.040 1.895 ;
        RECT  2.560 1.275 2.820 1.555 ;
        RECT  1.870 1.275 2.560 1.435 ;
        RECT  1.960 1.615 2.220 1.895 ;
        RECT  1.710 1.255 1.870 1.435 ;
        RECT  0.575 1.255 1.710 1.415 ;
        RECT  0.375 0.675 0.575 1.415 ;
        RECT  0.375 2.595 0.475 3.195 ;
        RECT  0.315 0.675 0.375 3.195 ;
        RECT  0.215 1.255 0.315 3.195 ;
    END
END NAND4BBX4

MACRO NAND4BBX2
    CLASS CORE ;
    FOREIGN NAND4BBX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.725 0.610 2.985 1.225 ;
        RECT  2.510 2.920 2.770 3.180 ;
        RECT  0.335 0.610 2.725 0.770 ;
        RECT  1.655 2.920 2.510 3.080 ;
        RECT  1.395 2.920 1.655 3.180 ;
        RECT  1.295 2.920 1.395 3.080 ;
        RECT  1.135 2.615 1.295 3.080 ;
        RECT  0.335 2.615 1.135 2.775 ;
        RECT  0.275 0.610 0.335 1.765 ;
        RECT  0.275 2.520 0.335 2.810 ;
        RECT  0.125 0.610 0.275 2.810 ;
        RECT  0.115 0.610 0.125 2.745 ;
        END
        ANTENNADIFFAREA     1.1755 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 2.520 4.015 2.810 ;
        RECT  2.525 2.525 3.805 2.685 ;
        RECT  2.365 2.525 2.525 2.740 ;
        RECT  1.635 2.580 2.365 2.740 ;
        RECT  1.475 2.105 1.635 2.740 ;
        RECT  1.315 1.705 1.475 2.265 ;
        END
        ANTENNAGATEAREA     0.3224 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.850 1.715 3.950 1.975 ;
        RECT  3.690 1.715 3.850 2.340 ;
        RECT  3.615 2.180 3.690 2.340 ;
        RECT  3.455 2.180 3.615 2.345 ;
        RECT  2.175 2.185 3.455 2.345 ;
        RECT  2.030 2.110 2.175 2.400 ;
        RECT  1.965 1.755 2.030 2.400 ;
        RECT  1.870 1.755 1.965 2.345 ;
        RECT  1.765 1.755 1.870 1.915 ;
        END
        ANTENNAGATEAREA     0.3224 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.725 1.760 4.935 2.400 ;
        RECT  4.635 1.760 4.725 2.270 ;
        RECT  4.535 1.760 4.635 2.020 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.795 1.930 ;
        RECT  0.535 1.670 0.585 1.930 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.425 -0.250 5.060 0.250 ;
        RECT  4.165 -0.250 4.425 1.135 ;
        RECT  1.490 -0.250 4.165 0.250 ;
        RECT  1.230 -0.250 1.490 0.405 ;
        RECT  0.000 -0.250 1.230 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.295 3.440 5.060 3.940 ;
        RECT  4.035 3.285 4.295 3.940 ;
        RECT  3.275 3.440 4.035 3.940 ;
        RECT  3.275 2.865 3.605 3.125 ;
        RECT  3.015 2.865 3.275 3.940 ;
        RECT  2.230 3.440 3.015 3.940 ;
        RECT  1.970 3.285 2.230 3.940 ;
        RECT  1.070 3.440 1.970 3.940 ;
        RECT  0.810 3.285 1.070 3.940 ;
        RECT  0.000 3.440 0.810 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.675 0.980 4.935 1.475 ;
        RECT  4.650 2.615 4.910 2.875 ;
        RECT  4.355 1.315 4.675 1.475 ;
        RECT  4.355 2.615 4.650 2.775 ;
        RECT  4.195 1.315 4.355 2.775 ;
        RECT  3.470 1.315 4.195 1.475 ;
        RECT  3.310 1.315 3.470 2.000 ;
        RECT  3.275 1.715 3.310 2.000 ;
        RECT  3.205 1.715 3.275 2.005 ;
        RECT  3.115 1.840 3.205 2.005 ;
        RECT  2.515 1.845 3.115 2.005 ;
        RECT  2.775 1.405 2.935 1.665 ;
        RECT  1.925 1.405 2.775 1.565 ;
        RECT  2.355 1.755 2.515 2.005 ;
        RECT  2.245 1.755 2.355 1.915 ;
        RECT  1.765 0.950 1.925 1.565 ;
        RECT  1.135 0.950 1.765 1.110 ;
        RECT  0.975 0.950 1.135 2.305 ;
        RECT  0.655 0.950 0.975 1.110 ;
        RECT  0.455 2.145 0.975 2.305 ;
    END
END NAND4BBX2

MACRO NAND4BBX1
    CLASS CORE ;
    FOREIGN NAND4BBX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.465 0.695 2.700 1.295 ;
        RECT  2.610 2.400 2.635 2.810 ;
        RECT  2.525 2.280 2.610 2.810 ;
        RECT  2.465 1.970 2.525 2.810 ;
        RECT  2.425 0.695 2.465 2.810 ;
        RECT  2.305 1.135 2.425 2.570 ;
        RECT  2.265 1.970 2.305 2.570 ;
        RECT  1.395 2.290 2.265 2.450 ;
        RECT  1.135 2.290 1.395 2.550 ;
        END
        ANTENNADIFFAREA     0.7380 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.865 1.770 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.520 1.510 1.570 1.770 ;
        RECT  1.310 1.420 1.520 1.770 ;
        RECT  1.255 1.420 1.310 1.580 ;
        RECT  1.045 1.290 1.255 1.580 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.290 0.370 1.770 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.065 3.590 1.770 ;
        RECT  3.310 1.510 3.345 1.770 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.360 -0.250 3.680 0.250 ;
        RECT  3.100 -0.250 3.360 0.405 ;
        RECT  0.890 -0.250 3.100 0.250 ;
        RECT  0.630 -0.250 0.890 0.405 ;
        RECT  0.000 -0.250 0.630 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.075 3.440 3.680 3.940 ;
        RECT  2.815 2.895 3.075 3.940 ;
        RECT  1.945 3.440 2.815 3.940 ;
        RECT  1.685 2.895 1.945 3.940 ;
        RECT  0.855 3.440 1.685 3.940 ;
        RECT  0.595 2.895 0.855 3.940 ;
        RECT  0.000 3.440 0.595 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.295 1.970 3.555 2.230 ;
        RECT  3.070 1.970 3.295 2.130 ;
        RECT  3.070 1.035 3.160 1.295 ;
        RECT  2.910 1.035 3.070 2.130 ;
        RECT  2.645 1.510 2.910 1.770 ;
        RECT  1.950 1.590 2.050 1.850 ;
        RECT  1.790 0.930 1.950 2.110 ;
        RECT  0.385 0.930 1.790 1.090 ;
        RECT  0.385 1.950 1.790 2.110 ;
        RECT  0.125 0.820 0.385 1.090 ;
        RECT  0.225 1.950 0.385 2.460 ;
        RECT  0.125 2.200 0.225 2.460 ;
    END
END NAND4BBX1

MACRO NAND4BBXL
    CLASS CORE ;
    FOREIGN NAND4BBXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.240 0.625 2.400 0.885 ;
        RECT  2.175 0.625 2.240 2.395 ;
        RECT  2.080 0.625 2.175 2.585 ;
        RECT  1.920 2.100 2.080 3.055 ;
        RECT  1.130 2.895 1.920 3.055 ;
        RECT  0.870 2.895 1.130 3.155 ;
        END
        ANTENNADIFFAREA     0.4097 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.285 0.865 1.770 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.355 1.390 1.810 ;
        RECT  1.045 1.290 1.255 1.810 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.285 0.370 1.770 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 1.495 3.110 1.995 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 -0.250 3.220 0.250 ;
        RECT  2.650 -0.250 2.910 0.405 ;
        RECT  0.930 -0.250 2.650 0.250 ;
        RECT  0.670 -0.250 0.930 0.405 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.525 3.440 3.220 3.940 ;
        RECT  2.265 3.285 2.525 3.940 ;
        RECT  1.710 3.440 2.265 3.940 ;
        RECT  1.450 3.285 1.710 3.940 ;
        RECT  0.580 3.440 1.450 3.940 ;
        RECT  0.320 3.285 0.580 3.940 ;
        RECT  0.000 3.440 0.320 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.835 2.610 3.095 2.870 ;
        RECT  2.650 0.940 2.910 1.310 ;
        RECT  2.580 2.610 2.835 2.770 ;
        RECT  2.580 1.150 2.650 1.310 ;
        RECT  2.420 1.150 2.580 2.770 ;
        RECT  1.740 1.660 1.870 1.920 ;
        RECT  1.580 0.920 1.740 2.150 ;
        RECT  0.385 0.920 1.580 1.080 ;
        RECT  0.580 1.990 1.580 2.150 ;
        RECT  0.320 1.970 0.580 2.230 ;
        RECT  0.125 0.820 0.385 1.080 ;
    END
END NAND4BBXL

MACRO NAND4BX4
    CLASS CORE ;
    FOREIGN NAND4BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.435 0.990 7.695 3.095 ;
        RECT  6.590 0.990 7.435 1.250 ;
        RECT  1.305 2.835 7.435 3.095 ;
        RECT  6.165 0.865 6.590 1.250 ;
        RECT  5.855 0.865 6.165 1.125 ;
        RECT  5.705 0.695 5.855 1.125 ;
        RECT  5.445 0.475 5.705 1.125 ;
        RECT  3.800 0.865 5.445 1.125 ;
        RECT  3.540 0.475 3.800 1.125 ;
        RECT  2.440 0.475 3.540 0.735 ;
        END
        ANTENNADIFFAREA     2.4518 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.150 1.925 7.235 2.400 ;
        RECT  7.050 1.635 7.150 2.400 ;
        RECT  6.890 1.635 7.050 2.615 ;
        RECT  1.260 2.455 6.890 2.615 ;
        RECT  1.100 1.610 1.260 2.615 ;
        RECT  1.045 1.610 1.100 2.175 ;
        RECT  1.000 1.610 1.045 1.870 ;
        END
        ANTENNAGATEAREA     0.7046 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 1.615 6.665 1.875 ;
        RECT  6.405 1.615 6.565 2.275 ;
        RECT  1.740 2.115 6.405 2.275 ;
        RECT  1.580 1.630 1.740 2.275 ;
        RECT  1.505 1.630 1.580 1.990 ;
        RECT  1.480 1.630 1.505 1.890 ;
        END
        ANTENNAGATEAREA     0.7046 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.180 1.615 6.185 1.875 ;
        RECT  5.925 1.615 6.180 1.935 ;
        RECT  5.220 1.775 5.925 1.935 ;
        RECT  4.925 1.685 5.220 1.935 ;
        RECT  3.320 1.775 4.925 1.935 ;
        RECT  3.040 1.685 3.320 1.935 ;
        RECT  2.220 1.775 3.040 1.935 ;
        RECT  2.175 1.615 2.220 1.935 ;
        RECT  1.960 1.290 2.175 1.935 ;
        END
        ANTENNAGATEAREA     0.7046 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.730 1.925 0.795 2.400 ;
        RECT  0.570 1.610 0.730 2.400 ;
        END
        ANTENNAGATEAREA     0.2743 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.225 -0.250 7.820 0.250 ;
        RECT  6.965 -0.250 7.225 0.795 ;
        RECT  4.260 -0.250 6.965 0.250 ;
        RECT  4.000 -0.250 4.260 0.685 ;
        RECT  1.115 -0.250 4.000 0.250 ;
        RECT  0.855 -0.250 1.115 0.735 ;
        RECT  0.000 -0.250 0.855 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.500 3.440 7.820 3.940 ;
        RECT  7.240 3.285 7.500 3.940 ;
        RECT  6.415 3.440 7.240 3.940 ;
        RECT  6.155 3.285 6.415 3.940 ;
        RECT  5.285 3.440 6.155 3.940 ;
        RECT  4.685 3.285 5.285 3.940 ;
        RECT  3.575 3.440 4.685 3.940 ;
        RECT  2.975 3.285 3.575 3.940 ;
        RECT  2.110 3.440 2.975 3.940 ;
        RECT  1.850 3.285 2.110 3.940 ;
        RECT  1.015 3.440 1.850 3.940 ;
        RECT  0.755 2.955 1.015 3.940 ;
        RECT  0.000 3.440 0.755 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.440 1.305 5.700 1.565 ;
        RECT  2.820 1.305 5.440 1.465 ;
        RECT  2.720 1.305 2.820 1.565 ;
        RECT  2.560 0.945 2.720 1.565 ;
        RECT  0.475 0.945 2.560 1.105 ;
        RECT  0.375 0.675 0.475 1.275 ;
        RECT  0.375 2.615 0.475 3.215 ;
        RECT  0.215 0.675 0.375 3.215 ;
    END
END NAND4BX4

MACRO NAND4BX2
    CLASS CORE ;
    FOREIGN NAND4BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 1.290 4.015 3.080 ;
        RECT  3.095 1.290 3.760 1.450 ;
        RECT  2.405 2.920 3.760 3.080 ;
        RECT  2.980 1.105 3.095 1.450 ;
        RECT  2.820 0.950 2.980 1.450 ;
        RECT  2.565 0.950 2.820 1.110 ;
        RECT  2.305 0.850 2.565 1.110 ;
        RECT  2.145 2.920 2.405 3.195 ;
        RECT  1.325 2.920 2.145 3.080 ;
        RECT  1.065 2.920 1.325 3.195 ;
        END
        ANTENNADIFFAREA     1.1324 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 2.580 3.580 2.740 ;
        RECT  1.135 2.110 1.255 2.740 ;
        RECT  1.095 1.705 1.135 2.740 ;
        RECT  0.975 1.705 1.095 2.405 ;
        RECT  0.910 1.705 0.975 1.965 ;
        END
        ANTENNAGATEAREA     0.3224 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.545 1.925 3.555 2.175 ;
        RECT  3.445 1.725 3.545 2.175 ;
        RECT  3.285 1.725 3.445 2.365 ;
        RECT  1.715 2.205 3.285 2.365 ;
        RECT  1.600 2.110 1.715 2.400 ;
        RECT  1.505 1.705 1.600 2.400 ;
        RECT  1.440 1.705 1.505 2.365 ;
        RECT  1.390 1.705 1.440 1.965 ;
        END
        ANTENNAGATEAREA     0.3224 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.795 1.700 3.095 2.005 ;
        RECT  2.100 1.845 2.795 2.005 ;
        RECT  1.940 1.755 2.100 2.005 ;
        RECT  1.820 1.755 1.940 1.915 ;
        END
        ANTENNAGATEAREA     0.3224 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 2.335 0.795 2.810 ;
        RECT  0.565 1.635 0.725 2.810 ;
        RECT  0.430 1.635 0.565 1.895 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 -0.250 4.140 0.250 ;
        RECT  3.755 -0.250 4.015 1.025 ;
        RECT  1.010 -0.250 3.755 0.250 ;
        RECT  0.750 -0.250 1.010 0.795 ;
        RECT  0.000 -0.250 0.750 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.945 3.440 4.140 3.940 ;
        RECT  2.685 3.285 2.945 3.940 ;
        RECT  1.865 3.440 2.685 3.940 ;
        RECT  1.605 3.285 1.865 3.940 ;
        RECT  0.785 3.440 1.605 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.305 1.295 2.565 1.665 ;
        RECT  0.470 1.295 2.305 1.455 ;
        RECT  0.250 1.010 0.470 1.455 ;
        RECT  0.250 2.075 0.385 2.675 ;
        RECT  0.210 1.010 0.250 2.675 ;
        RECT  0.125 1.295 0.210 2.675 ;
        RECT  0.090 1.295 0.125 2.235 ;
    END
END NAND4BX2

MACRO NAND4BX1
    CLASS CORE ;
    FOREIGN NAND4BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.695 2.635 2.585 ;
        RECT  2.585 0.695 2.610 2.730 ;
        RECT  2.425 0.480 2.585 2.730 ;
        RECT  2.235 2.570 2.425 2.730 ;
        RECT  1.975 2.570 2.235 2.830 ;
        RECT  1.295 2.670 1.975 2.830 ;
        RECT  1.135 2.670 1.295 3.230 ;
        RECT  1.035 3.070 1.135 3.230 ;
        END
        ANTENNADIFFAREA     0.9900 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.300 1.080 1.460 ;
        RECT  0.585 1.300 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.670 1.435 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.745 1.290 1.905 1.990 ;
        RECT  1.715 1.290 1.745 1.450 ;
        RECT  1.510 0.880 1.715 1.450 ;
        RECT  1.505 0.880 1.510 1.170 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.145 1.290 0.405 1.825 ;
        RECT  0.125 1.290 0.145 1.765 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 -0.250 2.760 0.250 ;
        RECT  0.660 -0.250 0.920 0.405 ;
        RECT  0.000 -0.250 0.660 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 3.440 2.760 3.940 ;
        RECT  2.375 3.285 2.635 3.940 ;
        RECT  1.835 3.440 2.375 3.940 ;
        RECT  1.575 3.285 1.835 3.940 ;
        RECT  0.405 3.440 1.575 3.940 ;
        RECT  0.145 3.285 0.405 3.940 ;
        RECT  0.000 3.440 0.145 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.085 0.535 2.245 2.390 ;
        RECT  1.260 0.535 2.085 0.695 ;
        RECT  0.385 2.230 2.085 2.390 ;
        RECT  1.100 0.535 1.260 1.010 ;
        RECT  0.385 0.850 1.100 1.010 ;
        RECT  0.125 0.850 0.385 1.110 ;
        RECT  0.225 2.230 0.385 2.920 ;
        RECT  0.125 2.660 0.225 2.920 ;
    END
END NAND4BX1

MACRO NAND4BXL
    CLASS CORE ;
    FOREIGN NAND4BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.480 0.825 2.640 2.875 ;
        RECT  2.425 0.825 2.480 1.170 ;
        RECT  2.230 2.715 2.480 2.875 ;
        RECT  2.375 0.825 2.425 1.085 ;
        RECT  1.970 2.610 2.230 2.875 ;
        RECT  1.255 2.715 1.970 2.875 ;
        RECT  0.995 2.715 1.255 3.090 ;
        END
        ANTENNADIFFAREA     0.5715 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.395 0.865 1.990 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.760 1.385 2.020 ;
        RECT  1.095 1.290 1.255 2.020 ;
        RECT  1.045 1.290 1.095 1.765 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.780 1.690 1.960 1.950 ;
        RECT  1.715 1.355 1.780 1.950 ;
        RECT  1.620 1.290 1.715 1.950 ;
        RECT  1.505 1.290 1.620 1.580 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.270 0.355 1.530 ;
        RECT  0.175 1.270 0.335 1.990 ;
        RECT  0.125 1.515 0.175 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.020 -0.250 2.760 0.250 ;
        RECT  0.760 -0.250 1.020 0.745 ;
        RECT  0.000 -0.250 0.760 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 3.440 2.760 3.940 ;
        RECT  2.375 3.285 2.635 3.940 ;
        RECT  1.805 3.440 2.375 3.940 ;
        RECT  1.545 3.285 1.805 3.940 ;
        RECT  0.745 3.440 1.545 3.940 ;
        RECT  0.485 3.285 0.745 3.940 ;
        RECT  0.000 3.440 0.485 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.140 1.350 2.300 2.430 ;
        RECT  2.120 1.350 2.140 1.510 ;
        RECT  0.385 2.270 2.140 2.430 ;
        RECT  1.960 0.925 2.120 1.510 ;
        RECT  0.410 0.925 1.960 1.085 ;
        RECT  0.150 0.825 0.410 1.085 ;
        RECT  0.225 2.270 0.385 2.975 ;
        RECT  0.125 2.715 0.225 2.975 ;
    END
END NAND4BXL

MACRO NAND3BX4
    CLASS CORE ;
    FOREIGN NAND3BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.910 0.585 4.935 2.335 ;
        RECT  4.650 0.585 4.910 2.465 ;
        RECT  4.380 0.585 4.650 1.205 ;
        RECT  4.475 2.110 4.650 2.465 ;
        RECT  4.450 2.110 4.475 2.585 ;
        RECT  4.365 2.225 4.450 2.585 ;
        RECT  2.235 0.585 4.380 0.825 ;
        RECT  4.105 2.225 4.365 3.185 ;
        RECT  3.055 2.535 4.105 2.735 ;
        RECT  2.455 2.535 3.055 2.795 ;
        RECT  1.405 2.535 2.455 2.735 ;
        RECT  1.975 0.555 2.235 0.825 ;
        RECT  1.145 2.535 1.405 3.135 ;
        END
        ANTENNADIFFAREA     2.7656 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 1.755 3.480 2.015 ;
        RECT  3.220 1.755 3.380 2.355 ;
        RECT  1.265 2.195 3.220 2.355 ;
        RECT  1.255 1.465 1.265 2.355 ;
        RECT  1.105 1.290 1.255 2.355 ;
        RECT  1.070 1.290 1.105 1.765 ;
        RECT  1.045 1.290 1.070 1.725 ;
        RECT  1.005 1.465 1.045 1.725 ;
        END
        ANTENNAGATEAREA     0.5954 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.825 1.755 3.960 2.015 ;
        RECT  3.665 1.415 3.825 2.015 ;
        RECT  2.885 1.415 3.665 1.575 ;
        RECT  2.725 1.415 2.885 2.015 ;
        RECT  2.625 1.725 2.725 2.015 ;
        RECT  1.745 1.855 2.625 2.015 ;
        RECT  1.715 1.755 1.745 2.015 ;
        RECT  1.505 1.700 1.715 2.015 ;
        RECT  1.485 1.755 1.505 2.015 ;
        END
        ANTENNAGATEAREA     0.5954 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 1.290 0.795 1.765 ;
        RECT  0.565 1.290 0.725 1.965 ;
        RECT  0.465 1.705 0.565 1.965 ;
        END
        ANTENNAGATEAREA     0.2522 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 -0.250 5.060 0.250 ;
        RECT  3.135 -0.250 3.395 0.405 ;
        RECT  1.065 -0.250 3.135 0.250 ;
        RECT  0.805 -0.250 1.065 0.745 ;
        RECT  0.000 -0.250 0.805 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.905 3.440 5.060 3.940 ;
        RECT  4.645 2.895 4.905 3.940 ;
        RECT  3.825 3.440 4.645 3.940 ;
        RECT  3.565 2.945 3.825 3.940 ;
        RECT  1.945 3.440 3.565 3.940 ;
        RECT  1.685 2.945 1.945 3.940 ;
        RECT  0.895 3.440 1.685 3.940 ;
        RECT  0.635 2.265 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.180 1.415 4.440 1.675 ;
        RECT  4.170 1.415 4.180 1.575 ;
        RECT  4.010 1.035 4.170 1.575 ;
        RECT  2.405 1.035 4.010 1.195 ;
        RECT  2.145 1.035 2.405 1.675 ;
        RECT  1.795 1.035 2.145 1.195 ;
        RECT  1.635 0.935 1.795 1.195 ;
        RECT  0.495 0.935 1.635 1.095 ;
        RECT  0.285 0.475 0.495 1.095 ;
        RECT  0.285 2.150 0.385 3.090 ;
        RECT  0.125 0.475 0.285 3.090 ;
    END
END NAND3BX4

MACRO NAND3BX2
    CLASS CORE ;
    FOREIGN NAND3BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.195 2.200 2.455 2.460 ;
        RECT  1.325 2.300 2.195 2.460 ;
        RECT  1.785 0.925 1.945 1.185 ;
        RECT  1.325 1.025 1.785 1.185 ;
        RECT  1.165 1.025 1.325 2.460 ;
        RECT  1.045 2.110 1.165 2.460 ;
        END
        ANTENNADIFFAREA     1.0504 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 2.205 2.995 2.465 ;
        RECT  2.735 2.205 2.895 2.835 ;
        RECT  0.865 2.675 2.735 2.835 ;
        RECT  0.865 1.405 0.985 1.665 ;
        RECT  0.705 1.405 0.865 2.835 ;
        RECT  0.585 1.925 0.705 2.400 ;
        END
        ANTENNAGATEAREA     0.2938 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 0.880 3.095 1.170 ;
        RECT  2.635 1.010 2.885 1.170 ;
        RECT  2.475 1.010 2.635 2.015 ;
        RECT  1.665 1.855 2.475 2.015 ;
        RECT  1.505 1.725 1.665 2.015 ;
        END
        ANTENNAGATEAREA     0.2938 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.800 0.525 3.060 ;
        RECT  0.125 2.800 0.335 3.220 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.220 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.785 -0.250 2.835 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 3.440 3.220 3.940 ;
        RECT  1.655 3.285 1.915 3.940 ;
        RECT  0.825 3.440 1.655 3.940 ;
        RECT  0.565 3.285 0.825 3.940 ;
        RECT  0.000 3.440 0.565 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.135 0.585 2.295 1.675 ;
        RECT  0.385 0.585 2.135 0.745 ;
        RECT  1.935 1.415 2.135 1.675 ;
        RECT  0.225 0.585 0.385 2.505 ;
        RECT  0.125 1.035 0.225 1.295 ;
        RECT  0.125 2.245 0.225 2.505 ;
    END
END NAND3BX2

MACRO NAND3BX1
    CLASS CORE ;
    FOREIGN NAND3BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 0.825 2.210 1.765 ;
        RECT  2.090 0.825 2.175 3.145 ;
        RECT  2.050 0.725 2.090 3.145 ;
        RECT  1.830 0.725 2.050 0.985 ;
        RECT  1.965 1.605 2.050 3.145 ;
        RECT  1.915 2.885 1.965 3.145 ;
        RECT  1.300 2.885 1.915 3.045 ;
        RECT  1.040 2.855 1.300 3.115 ;
        END
        ANTENNADIFFAREA     0.7749 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.075 2.110 1.255 2.400 ;
        RECT  0.915 1.505 1.075 2.400 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.665 1.925 1.715 2.400 ;
        RECT  1.505 1.645 1.665 2.400 ;
        RECT  1.425 1.645 1.505 1.905 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.570 1.545 0.730 2.680 ;
        RECT  0.430 1.545 0.570 1.805 ;
        RECT  0.335 2.520 0.570 2.680 ;
        RECT  0.125 2.520 0.335 2.810 ;
        END
        ANTENNAGATEAREA     0.0650 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.925 -0.250 2.300 0.250 ;
        RECT  0.665 -0.250 0.925 0.405 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 3.440 2.300 3.940 ;
        RECT  0.525 2.895 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.710 1.165 1.870 1.425 ;
        RECT  1.620 1.165 1.710 1.325 ;
        RECT  1.460 0.895 1.620 1.325 ;
        RECT  0.440 0.895 1.460 1.055 ;
        RECT  0.340 0.795 0.440 1.055 ;
        RECT  0.250 1.985 0.385 2.275 ;
        RECT  0.250 0.795 0.340 1.365 ;
        RECT  0.180 0.795 0.250 2.275 ;
        RECT  0.125 1.205 0.180 2.275 ;
        RECT  0.090 1.205 0.125 2.145 ;
    END
END NAND3BX1

MACRO NAND3BXL
    CLASS CORE ;
    FOREIGN NAND3BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.900 2.175 2.810 ;
        RECT  2.015 0.900 2.150 2.985 ;
        RECT  1.915 0.900 2.015 1.060 ;
        RECT  1.965 1.925 2.015 2.985 ;
        RECT  1.870 2.725 1.965 2.985 ;
        RECT  0.995 2.775 1.870 2.935 ;
        END
        ANTENNADIFFAREA     0.5881 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.860 1.415 1.020 2.590 ;
        RECT  0.795 2.430 0.860 2.590 ;
        RECT  0.585 2.430 0.795 2.810 ;
        END
        ANTENNAGATEAREA     0.0897 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.110 1.715 2.400 ;
        RECT  1.500 2.110 1.505 2.270 ;
        RECT  1.340 1.735 1.500 2.270 ;
        END
        ANTENNAGATEAREA     0.0897 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.090 0.335 1.895 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 -0.250 2.300 0.250 ;
        RECT  0.640 -0.250 0.900 0.405 ;
        RECT  0.000 -0.250 0.640 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.615 3.440 2.300 3.940 ;
        RECT  0.635 3.285 1.615 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.650 1.240 1.810 1.500 ;
        RECT  1.590 1.240 1.650 1.400 ;
        RECT  1.430 0.900 1.590 1.400 ;
        RECT  0.680 0.900 1.430 1.060 ;
        RECT  0.520 0.635 0.680 2.245 ;
        RECT  0.385 0.635 0.520 0.855 ;
        RECT  0.285 2.085 0.520 2.245 ;
        RECT  0.125 0.595 0.385 0.855 ;
        RECT  0.285 3.055 0.385 3.215 ;
        RECT  0.125 2.085 0.285 3.215 ;
    END
END NAND3BXL

MACRO NAND2BX4
    CLASS CORE ;
    FOREIGN NAND2BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.545 0.880 3.555 2.175 ;
        RECT  3.370 0.880 3.545 2.395 ;
        RECT  3.345 0.665 3.370 2.395 ;
        RECT  3.095 0.665 3.345 1.265 ;
        RECT  2.425 2.195 3.345 2.395 ;
        RECT  3.070 0.665 3.095 1.195 ;
        RECT  1.715 0.995 3.070 1.195 ;
        RECT  2.165 2.195 2.425 3.160 ;
        RECT  1.405 2.195 2.165 2.395 ;
        RECT  1.455 0.555 1.715 1.195 ;
        RECT  1.145 2.195 1.405 3.160 ;
        END
        ANTENNADIFFAREA     1.4444 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.305 1.375 2.565 1.635 ;
        RECT  1.255 1.375 2.305 1.535 ;
        RECT  1.065 1.290 1.255 1.580 ;
        RECT  0.855 1.290 1.065 1.635 ;
        END
        ANTENNAGATEAREA     0.6019 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.445 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2431 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.535 -0.250 4.140 0.250 ;
        RECT  2.275 -0.250 2.535 0.815 ;
        RECT  0.895 -0.250 2.275 0.250 ;
        RECT  0.635 -0.250 0.895 0.825 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 3.440 4.140 3.940 ;
        RECT  2.675 2.590 2.935 3.940 ;
        RECT  1.915 3.440 2.675 3.940 ;
        RECT  1.655 2.590 1.915 3.940 ;
        RECT  0.895 3.440 1.655 3.940 ;
        RECT  0.635 2.535 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.975 1.675 3.135 1.975 ;
        RECT  1.745 1.815 2.975 1.975 ;
        RECT  1.485 1.725 1.745 1.975 ;
        RECT  0.675 1.815 1.485 1.975 ;
        RECT  0.515 1.005 0.675 2.330 ;
        RECT  0.385 1.005 0.515 1.265 ;
        RECT  0.385 2.170 0.515 2.330 ;
        RECT  0.125 0.665 0.385 1.265 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END NAND2BX4

MACRO NAND2BX2
    CLASS CORE ;
    FOREIGN NAND2BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.515 2.635 2.175 ;
        RECT  2.425 1.250 2.585 2.355 ;
        RECT  2.165 1.250 2.425 1.410 ;
        RECT  1.595 2.195 2.425 2.355 ;
        RECT  2.005 0.780 2.165 1.410 ;
        RECT  1.775 0.780 2.005 0.940 ;
        RECT  1.515 0.680 1.775 0.940 ;
        RECT  1.335 2.195 1.595 3.215 ;
        END
        ANTENNADIFFAREA     0.7228 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 1.595 2.245 1.990 ;
        RECT  1.255 1.830 1.985 1.990 ;
        RECT  1.220 1.700 1.255 1.990 ;
        RECT  0.960 1.595 1.220 1.990 ;
        END
        ANTENNAGATEAREA     0.3185 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.495 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1209 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.605 -0.250 2.760 0.250 ;
        RECT  2.345 -0.250 2.605 0.885 ;
        RECT  0.905 -0.250 2.345 0.250 ;
        RECT  0.905 0.630 0.940 0.890 ;
        RECT  0.645 -0.250 0.905 0.890 ;
        RECT  0.000 -0.250 0.645 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.135 3.440 2.760 3.940 ;
        RECT  1.875 2.545 2.135 3.940 ;
        RECT  1.050 3.440 1.875 3.940 ;
        RECT  0.790 2.550 1.050 3.940 ;
        RECT  0.000 3.440 0.790 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.600 1.310 1.730 1.570 ;
        RECT  1.440 1.120 1.600 1.570 ;
        RECT  0.780 1.120 1.440 1.280 ;
        RECT  0.620 1.120 0.780 2.370 ;
        RECT  0.385 1.120 0.620 1.280 ;
        RECT  0.385 2.210 0.620 2.370 ;
        RECT  0.125 0.995 0.385 1.280 ;
        RECT  0.125 2.210 0.385 2.625 ;
    END
END NAND2BX2

MACRO NAND2BX1
    CLASS CORE ;
    FOREIGN NAND2BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 0.880 1.725 2.630 ;
        RECT  1.505 0.880 1.565 1.355 ;
        RECT  1.530 2.335 1.565 2.630 ;
        RECT  1.295 2.470 1.530 2.630 ;
        RECT  1.455 0.880 1.505 1.160 ;
        RECT  1.035 2.470 1.295 2.730 ;
        END
        ANTENNADIFFAREA     0.4404 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.780 1.790 0.925 1.950 ;
        RECT  0.780 1.290 0.795 1.580 ;
        RECT  0.620 1.290 0.780 1.950 ;
        RECT  0.585 1.290 0.620 1.580 ;
        END
        ANTENNAGATEAREA     0.1586 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.510 0.385 1.770 ;
        RECT  0.125 1.510 0.335 2.215 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.805 -0.250 1.840 0.250 ;
        RECT  0.545 -0.250 0.805 0.745 ;
        RECT  0.000 -0.250 0.545 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.695 3.440 1.840 3.940 ;
        RECT  1.435 3.285 1.695 3.940 ;
        RECT  0.960 3.440 1.435 3.940 ;
        RECT  0.700 3.235 0.960 3.940 ;
        RECT  0.000 3.440 0.700 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.265 1.750 1.385 2.010 ;
        RECT  1.105 0.930 1.265 2.290 ;
        RECT  0.385 0.930 1.105 1.090 ;
        RECT  0.685 2.130 1.105 2.290 ;
        RECT  0.525 2.130 0.685 2.585 ;
        RECT  0.385 2.425 0.525 2.585 ;
        RECT  0.125 0.930 0.385 1.295 ;
        RECT  0.225 2.425 0.385 3.080 ;
        RECT  0.125 2.820 0.225 3.080 ;
    END
END NAND2BX1

MACRO NAND2BXL
    CLASS CORE ;
    FOREIGN NAND2BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 0.480 1.715 2.810 ;
        RECT  1.500 0.480 1.555 1.325 ;
        RECT  1.505 1.950 1.555 2.810 ;
        RECT  1.400 2.620 1.505 2.810 ;
        RECT  1.455 0.480 1.500 0.740 ;
        RECT  1.140 2.620 1.400 2.880 ;
        END
        ANTENNADIFFAREA     0.5012 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.600 0.930 1.860 ;
        RECT  0.635 1.290 0.795 1.860 ;
        RECT  0.585 1.290 0.635 1.765 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.325 0.375 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 -0.250 1.840 0.250 ;
        RECT  0.660 -0.250 0.920 0.405 ;
        RECT  0.000 -0.250 0.660 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.395 3.440 1.840 3.940 ;
        RECT  1.135 3.285 1.395 3.940 ;
        RECT  0.815 3.440 1.135 3.940 ;
        RECT  0.555 2.895 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.270 1.505 1.360 1.765 ;
        RECT  1.110 0.680 1.270 2.340 ;
        RECT  0.410 0.680 1.110 0.840 ;
        RECT  0.900 2.180 1.110 2.340 ;
        RECT  0.740 2.180 0.900 2.450 ;
        RECT  0.385 2.290 0.740 2.450 ;
        RECT  0.250 0.430 0.410 0.840 ;
        RECT  0.125 2.290 0.385 2.550 ;
        RECT  0.150 0.430 0.250 0.590 ;
    END
END NAND2BXL

MACRO NAND4X8
    CLASS CORE ;
    FOREIGN NAND4X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.065 1.515 14.135 3.095 ;
        RECT  13.655 1.180 14.065 3.095 ;
        RECT  13.215 1.180 13.655 1.580 ;
        RECT  2.150 2.805 13.655 3.095 ;
        RECT  12.805 0.880 13.215 1.580 ;
        RECT  12.545 0.545 12.805 1.580 ;
        RECT  11.335 0.545 12.545 0.805 ;
        RECT  7.345 0.585 11.335 0.805 ;
        RECT  7.085 0.585 7.345 1.185 ;
        RECT  7.025 0.695 7.085 1.185 ;
        RECT  4.235 0.875 7.025 1.185 ;
        RECT  3.975 0.585 4.235 1.185 ;
        RECT  2.090 2.745 2.150 3.095 ;
        RECT  2.075 2.250 2.090 3.095 ;
        RECT  1.800 2.250 2.075 3.190 ;
        RECT  1.010 2.250 1.800 2.540 ;
        RECT  0.720 2.250 1.010 3.190 ;
        RECT  0.365 2.250 0.720 2.590 ;
        RECT  0.365 0.615 0.465 1.215 ;
        RECT  0.205 0.615 0.365 2.590 ;
        RECT  0.125 1.105 0.205 2.175 ;
        END
        ANTENNADIFFAREA     5.2094 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.065 2.255 13.325 2.615 ;
        RECT  9.535 2.455 13.065 2.615 ;
        RECT  9.275 2.320 9.535 2.615 ;
        RECT  2.635 2.455 9.275 2.615 ;
        RECT  2.475 1.705 2.635 2.615 ;
        RECT  2.425 1.705 2.475 2.400 ;
        RECT  2.375 1.705 2.425 1.965 ;
        END
        ANTENNAGATEAREA     1.3494 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.585 2.015 12.845 2.275 ;
        RECT  10.485 2.115 12.585 2.275 ;
        RECT  10.325 1.750 10.485 2.275 ;
        RECT  10.215 1.750 10.325 1.915 ;
        RECT  8.400 1.755 10.215 1.915 ;
        RECT  8.240 1.755 8.400 2.275 ;
        RECT  3.115 2.115 8.240 2.275 ;
        RECT  2.955 1.365 3.115 2.275 ;
        RECT  2.885 1.365 2.955 1.765 ;
        RECT  2.855 1.365 2.885 1.645 ;
        RECT  2.175 1.365 2.855 1.525 ;
        RECT  2.125 1.290 2.175 1.765 ;
        RECT  1.965 1.290 2.125 1.865 ;
        RECT  1.785 1.705 1.965 1.865 ;
        RECT  1.525 1.705 1.785 1.965 ;
        END
        ANTENNAGATEAREA     1.3494 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.845 1.755 12.365 1.915 ;
        RECT  10.685 1.365 10.845 1.915 ;
        RECT  8.050 1.365 10.685 1.525 ;
        RECT  7.890 1.365 8.050 1.935 ;
        RECT  7.760 1.755 7.890 1.935 ;
        RECT  6.865 1.775 7.760 1.935 ;
        RECT  6.655 1.755 6.865 1.935 ;
        RECT  5.530 1.755 6.655 1.915 ;
        RECT  4.625 1.755 5.530 1.935 ;
        RECT  3.595 1.775 4.625 1.935 ;
        RECT  3.455 1.755 3.595 1.935 ;
        RECT  3.295 0.930 3.455 1.935 ;
        RECT  1.300 0.930 3.295 1.090 ;
        RECT  1.140 0.930 1.300 1.645 ;
        RECT  1.045 1.290 1.140 1.645 ;
        RECT  1.040 1.385 1.045 1.645 ;
        END
        ANTENNAGATEAREA     1.3494 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.690 1.205 11.790 1.465 ;
        RECT  11.530 1.015 11.690 1.465 ;
        RECT  7.705 1.015 11.530 1.175 ;
        RECT  7.545 1.015 7.705 1.575 ;
        RECT  7.515 1.415 7.545 1.575 ;
        RECT  7.255 1.415 7.515 1.595 ;
        RECT  4.405 1.415 7.255 1.575 ;
        RECT  4.145 1.415 4.405 1.595 ;
        RECT  3.795 1.415 4.145 1.575 ;
        RECT  3.635 0.590 3.795 1.575 ;
        RECT  0.860 0.590 3.635 0.750 ;
        RECT  0.795 0.590 0.860 1.645 ;
        RECT  0.700 0.590 0.795 1.990 ;
        RECT  0.600 1.435 0.700 1.990 ;
        RECT  0.585 1.700 0.600 1.990 ;
        END
        ANTENNAGATEAREA     1.3494 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.750 -0.250 14.260 0.250 ;
        RECT  13.490 -0.250 13.750 0.880 ;
        RECT  13.275 -0.250 13.490 0.405 ;
        RECT  9.700 -0.250 13.275 0.250 ;
        RECT  9.440 -0.250 9.700 0.405 ;
        RECT  9.010 -0.250 9.440 0.250 ;
        RECT  8.750 -0.250 9.010 0.405 ;
        RECT  5.875 -0.250 8.750 0.250 ;
        RECT  5.615 -0.250 5.875 0.405 ;
        RECT  2.435 -0.250 5.615 0.250 ;
        RECT  2.175 -0.250 2.435 0.405 ;
        RECT  0.000 -0.250 2.175 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.925 3.440 14.260 3.940 ;
        RECT  11.665 3.285 11.925 3.940 ;
        RECT  10.845 3.440 11.665 3.940 ;
        RECT  10.585 3.285 10.845 3.940 ;
        RECT  9.740 3.440 10.585 3.940 ;
        RECT  9.140 3.285 9.740 3.940 ;
        RECT  8.225 3.440 9.140 3.940 ;
        RECT  7.965 3.285 8.225 3.940 ;
        RECT  7.120 3.440 7.965 3.940 ;
        RECT  6.860 3.285 7.120 3.940 ;
        RECT  4.800 3.440 6.860 3.940 ;
        RECT  4.540 3.285 4.800 3.940 ;
        RECT  3.695 3.440 4.540 3.940 ;
        RECT  3.435 3.285 3.695 3.940 ;
        RECT  2.615 3.440 3.435 3.940 ;
        RECT  2.355 3.285 2.615 3.940 ;
        RECT  1.535 3.440 2.355 3.940 ;
        RECT  1.275 2.820 1.535 3.940 ;
        RECT  0.410 3.440 1.275 3.940 ;
        RECT  0.150 2.820 0.410 3.940 ;
        RECT  0.000 3.440 0.150 3.940 ;
        END
    END VDD
END NAND4X8

MACRO NAND4X6
    CLASS CORE ;
    FOREIGN NAND4X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.530 0.875 9.535 2.585 ;
        RECT  9.240 0.875 9.530 3.095 ;
        RECT  8.865 0.875 9.240 1.580 ;
        RECT  2.150 2.805 9.240 3.095 ;
        RECT  7.345 0.875 8.865 1.185 ;
        RECT  7.085 0.585 7.345 1.185 ;
        RECT  7.025 0.695 7.085 1.185 ;
        RECT  4.235 0.875 7.025 1.185 ;
        RECT  3.975 0.585 4.235 1.185 ;
        RECT  2.090 2.745 2.150 3.095 ;
        RECT  2.075 2.215 2.090 3.095 ;
        RECT  1.800 2.215 2.075 3.195 ;
        RECT  1.080 2.215 1.800 2.505 ;
        RECT  0.770 2.215 1.080 3.195 ;
        RECT  0.420 2.215 0.770 2.505 ;
        RECT  0.420 0.950 0.465 1.250 ;
        RECT  0.130 0.950 0.420 2.505 ;
        RECT  0.125 1.105 0.130 2.505 ;
        END
        ANTENNADIFFAREA     3.6283 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.890 1.765 9.050 2.615 ;
        RECT  2.635 2.455 8.890 2.615 ;
        RECT  2.475 1.705 2.635 2.615 ;
        RECT  2.425 1.705 2.475 2.400 ;
        RECT  2.375 1.705 2.425 1.965 ;
        END
        ANTENNAGATEAREA     0.9776 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.400 1.765 8.500 2.025 ;
        RECT  8.240 1.765 8.400 2.275 ;
        RECT  3.115 2.115 8.240 2.275 ;
        RECT  2.955 1.365 3.115 2.275 ;
        RECT  2.885 1.365 2.955 1.765 ;
        RECT  2.855 1.365 2.885 1.645 ;
        RECT  2.175 1.365 2.855 1.525 ;
        RECT  2.125 1.290 2.175 1.765 ;
        RECT  1.965 1.290 2.125 1.865 ;
        RECT  1.785 1.705 1.965 1.865 ;
        RECT  1.525 1.705 1.785 1.965 ;
        END
        ANTENNAGATEAREA     0.9776 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 1.775 8.020 1.935 ;
        RECT  4.625 1.755 4.885 1.935 ;
        RECT  3.595 1.775 4.625 1.935 ;
        RECT  3.455 1.755 3.595 1.935 ;
        RECT  3.295 0.930 3.455 1.935 ;
        RECT  1.300 0.930 3.295 1.090 ;
        RECT  1.140 0.930 1.300 1.645 ;
        RECT  1.045 1.290 1.140 1.645 ;
        RECT  1.040 1.385 1.045 1.645 ;
        END
        ANTENNAGATEAREA     0.9776 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.255 1.415 7.515 1.595 ;
        RECT  4.405 1.415 7.255 1.575 ;
        RECT  4.145 1.415 4.405 1.595 ;
        RECT  3.795 1.415 4.145 1.575 ;
        RECT  3.635 0.590 3.795 1.575 ;
        RECT  0.860 0.590 3.635 0.750 ;
        RECT  0.795 0.590 0.860 1.960 ;
        RECT  0.700 0.470 0.795 1.960 ;
        RECT  0.585 0.470 0.700 0.760 ;
        RECT  0.610 1.700 0.700 1.960 ;
        END
        ANTENNAGATEAREA     0.9776 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.010 -0.250 9.660 0.250 ;
        RECT  8.750 -0.250 9.010 0.405 ;
        RECT  5.875 -0.250 8.750 0.250 ;
        RECT  5.615 -0.250 5.875 0.405 ;
        RECT  2.435 -0.250 5.615 0.250 ;
        RECT  2.175 -0.250 2.435 0.405 ;
        RECT  0.000 -0.250 2.175 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.470 3.440 9.660 3.940 ;
        RECT  9.210 3.285 9.470 3.940 ;
        RECT  8.390 3.440 9.210 3.940 ;
        RECT  8.130 3.285 8.390 3.940 ;
        RECT  7.285 3.440 8.130 3.940 ;
        RECT  7.025 3.285 7.285 3.940 ;
        RECT  4.800 3.440 7.025 3.940 ;
        RECT  4.540 3.285 4.800 3.940 ;
        RECT  3.695 3.440 4.540 3.940 ;
        RECT  3.435 3.285 3.695 3.940 ;
        RECT  2.615 3.440 3.435 3.940 ;
        RECT  2.355 3.285 2.615 3.940 ;
        RECT  1.565 3.440 2.355 3.940 ;
        RECT  1.305 2.935 1.565 3.940 ;
        RECT  0.470 3.440 1.305 3.940 ;
        RECT  0.210 2.890 0.470 3.940 ;
        RECT  0.000 3.440 0.210 3.940 ;
        END
    END VDD
END NAND4X6

MACRO NAND4X4
    CLASS CORE ;
    FOREIGN NAND4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.975 1.085 7.235 3.095 ;
        RECT  5.670 1.085 6.975 1.325 ;
        RECT  0.635 2.835 6.975 3.095 ;
        RECT  5.240 0.925 5.670 1.325 ;
        RECT  5.215 0.925 5.240 1.165 ;
        RECT  5.035 0.880 5.215 1.165 ;
        RECT  4.775 0.550 5.035 1.165 ;
        RECT  4.725 0.695 4.775 1.165 ;
        RECT  3.120 0.925 4.725 1.165 ;
        RECT  2.880 0.870 3.120 1.165 ;
        RECT  2.175 0.870 2.880 1.110 ;
        RECT  2.150 0.695 2.175 1.110 ;
        RECT  1.890 0.510 2.150 1.110 ;
        END
        ANTENNADIFFAREA     2.4503 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.380 1.510 6.480 1.770 ;
        RECT  6.220 1.510 6.380 2.630 ;
        RECT  6.105 2.335 6.220 2.630 ;
        RECT  3.590 2.470 6.105 2.630 ;
        RECT  3.330 2.410 3.590 2.630 ;
        RECT  0.405 2.470 3.330 2.630 ;
        RECT  0.245 1.635 0.405 2.630 ;
        RECT  0.145 1.635 0.245 2.400 ;
        RECT  0.125 1.890 0.145 2.400 ;
        END
        ANTENNAGATEAREA     0.7046 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.895 1.615 5.995 1.875 ;
        RECT  5.735 1.615 5.895 2.290 ;
        RECT  4.070 2.130 5.735 2.290 ;
        RECT  3.810 2.025 4.070 2.290 ;
        RECT  3.110 2.025 3.810 2.185 ;
        RECT  2.850 2.025 3.110 2.275 ;
        RECT  1.190 2.115 2.850 2.275 ;
        RECT  1.030 1.615 1.190 2.275 ;
        RECT  0.930 1.615 1.030 1.990 ;
        RECT  0.585 1.700 0.930 1.990 ;
        END
        ANTENNAGATEAREA     0.7046 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.255 1.615 5.515 1.950 ;
        RECT  4.550 1.790 5.255 1.950 ;
        RECT  4.255 1.685 4.550 1.950 ;
        RECT  2.650 1.685 4.255 1.845 ;
        RECT  2.370 1.685 2.650 1.935 ;
        RECT  1.670 1.775 2.370 1.935 ;
        RECT  1.570 1.615 1.670 1.935 ;
        RECT  1.410 1.010 1.570 1.935 ;
        RECT  1.255 1.010 1.410 1.170 ;
        RECT  1.045 0.880 1.255 1.170 ;
        END
        ANTENNAGATEAREA     0.7046 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.770 1.345 5.030 1.610 ;
        RECT  2.175 1.345 4.770 1.505 ;
        RECT  1.965 1.290 2.175 1.580 ;
        RECT  1.890 1.315 1.965 1.575 ;
        END
        ANTENNAGATEAREA     0.7046 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.480 -0.250 7.360 0.250 ;
        RECT  6.220 -0.250 6.480 0.795 ;
        RECT  3.590 -0.250 6.220 0.250 ;
        RECT  3.330 -0.250 3.590 0.735 ;
        RECT  0.710 -0.250 3.330 0.250 ;
        RECT  0.450 -0.250 0.710 1.075 ;
        RECT  0.000 -0.250 0.450 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.830 3.440 7.360 3.940 ;
        RECT  6.570 3.285 6.830 3.940 ;
        RECT  5.745 3.440 6.570 3.940 ;
        RECT  5.485 3.285 5.745 3.940 ;
        RECT  4.660 3.440 5.485 3.940 ;
        RECT  4.060 3.285 4.660 3.940 ;
        RECT  2.860 3.440 4.060 3.940 ;
        RECT  2.260 3.285 2.860 3.940 ;
        RECT  1.440 3.440 2.260 3.940 ;
        RECT  1.180 3.285 1.440 3.940 ;
        RECT  0.385 3.440 1.180 3.940 ;
        RECT  0.125 2.935 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND4X4

MACRO NAND4X2
    CLASS CORE ;
    FOREIGN NAND4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 1.695 3.565 3.055 ;
        RECT  3.095 1.695 3.405 1.855 ;
        RECT  3.345 2.745 3.405 3.055 ;
        RECT  1.975 2.895 3.345 3.055 ;
        RECT  3.045 0.695 3.095 1.855 ;
        RECT  2.935 0.540 3.045 1.855 ;
        RECT  2.885 0.540 2.935 1.355 ;
        RECT  2.100 0.540 2.885 0.700 ;
        RECT  1.840 0.540 2.100 0.945 ;
        RECT  1.715 2.895 1.975 3.195 ;
        RECT  0.895 2.895 1.715 3.055 ;
        RECT  0.635 2.895 0.895 3.195 ;
        END
        ANTENNADIFFAREA     1.1134 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 2.035 3.225 2.295 ;
        RECT  2.965 2.035 3.125 2.665 ;
        RECT  2.885 2.335 2.965 2.665 ;
        RECT  0.405 2.505 2.885 2.665 ;
        RECT  0.245 1.465 0.405 2.665 ;
        RECT  0.125 1.465 0.245 2.175 ;
        END
        ANTENNAGATEAREA     0.3172 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.645 1.725 2.745 1.985 ;
        RECT  2.485 1.725 2.645 2.325 ;
        RECT  1.040 2.165 2.485 2.325 ;
        RECT  0.880 1.725 1.040 2.325 ;
        RECT  0.795 1.725 0.880 1.990 ;
        RECT  0.585 1.700 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.3172 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.450 1.725 1.635 1.985 ;
        RECT  1.290 1.010 1.450 1.985 ;
        RECT  1.255 1.010 1.290 1.170 ;
        RECT  1.045 0.880 1.255 1.170 ;
        END
        ANTENNAGATEAREA     0.3172 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.550 0.880 2.635 1.170 ;
        RECT  2.390 0.880 2.550 1.545 ;
        RECT  2.115 1.385 2.390 1.545 ;
        RECT  1.855 1.385 2.115 1.665 ;
        END
        ANTENNAGATEAREA     0.3172 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.545 -0.250 3.680 0.250 ;
        RECT  3.285 -0.250 3.545 1.285 ;
        RECT  0.540 -0.250 3.285 0.250 ;
        RECT  0.280 -0.250 0.540 1.285 ;
        RECT  0.000 -0.250 0.280 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 3.440 3.680 3.940 ;
        RECT  2.255 3.285 2.855 3.940 ;
        RECT  1.435 3.440 2.255 3.940 ;
        RECT  1.175 3.285 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.935 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND4X2

MACRO NAND4X1
    CLASS CORE ;
    FOREIGN NAND4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 0.965 2.205 1.905 ;
        RECT  2.045 0.525 2.175 2.400 ;
        RECT  1.915 0.525 2.045 1.125 ;
        RECT  2.015 1.745 2.045 2.400 ;
        RECT  1.965 2.110 2.015 2.400 ;
        RECT  1.775 2.185 1.965 2.395 ;
        RECT  1.505 2.185 1.775 2.785 ;
        RECT  0.795 2.185 1.505 2.345 ;
        RECT  0.525 2.185 0.795 2.785 ;
        END
        ANTENNADIFFAREA     0.9336 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.395 0.375 1.990 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.395 0.925 2.005 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.295 1.745 1.435 2.005 ;
        RECT  1.135 0.880 1.295 2.005 ;
        RECT  1.045 0.880 1.135 1.170 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.305 1.865 1.565 ;
        RECT  1.555 0.880 1.715 1.565 ;
        RECT  1.505 0.880 1.555 1.355 ;
        END
        ANTENNAGATEAREA     0.1794 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.250 2.300 0.250 ;
        RECT  0.125 -0.250 0.385 1.195 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 3.440 2.300 3.940 ;
        RECT  1.915 3.285 2.175 3.940 ;
        RECT  1.410 3.440 1.915 3.940 ;
        RECT  1.150 3.285 1.410 3.940 ;
        RECT  0.385 3.440 1.150 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND4X1

MACRO NAND4XL
    CLASS CORE ;
    FOREIGN NAND4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.030 0.935 2.190 2.585 ;
        RECT  1.965 0.935 2.030 1.580 ;
        RECT  1.990 2.335 2.030 2.585 ;
        RECT  1.775 2.425 1.990 2.585 ;
        RECT  1.915 0.935 1.965 1.195 ;
        RECT  1.515 2.425 1.775 2.720 ;
        RECT  0.785 2.425 1.515 2.585 ;
        RECT  0.525 2.425 0.785 2.720 ;
        END
        ANTENNADIFFAREA     0.5061 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.795 0.370 2.055 ;
        RECT  0.110 1.795 0.335 2.400 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.725 0.885 1.985 ;
        RECT  0.610 0.880 0.795 1.985 ;
        RECT  0.585 0.880 0.610 1.725 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.725 1.420 1.985 ;
        RECT  1.070 0.880 1.255 1.985 ;
        RECT  1.045 0.880 1.070 1.355 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.775 1.760 1.850 2.020 ;
        RECT  1.715 1.375 1.775 2.020 ;
        RECT  1.615 0.880 1.715 2.020 ;
        RECT  1.555 0.880 1.615 1.535 ;
        RECT  1.505 0.880 1.555 1.170 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.250 2.300 0.250 ;
        RECT  0.125 -0.250 0.385 1.135 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 3.440 2.300 3.940 ;
        RECT  1.915 3.285 2.175 3.940 ;
        RECT  1.440 3.440 1.915 3.940 ;
        RECT  1.180 3.285 1.440 3.940 ;
        RECT  0.385 3.440 1.180 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND4XL

MACRO NAND3X8
    CLASS CORE ;
    FOREIGN NAND3X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.715 1.180 9.075 3.100 ;
        RECT  8.675 1.180 8.715 3.040 ;
        RECT  8.615 1.180 8.675 1.580 ;
        RECT  8.590 2.520 8.675 3.040 ;
        RECT  7.945 0.585 8.615 1.580 ;
        RECT  7.970 2.655 8.590 3.040 ;
        RECT  7.895 2.595 7.970 3.040 ;
        RECT  3.135 0.585 7.945 0.985 ;
        RECT  7.635 2.595 7.895 3.195 ;
        RECT  6.815 2.655 7.635 3.025 ;
        RECT  6.555 2.595 6.815 3.195 ;
        RECT  5.735 2.655 6.555 3.025 ;
        RECT  5.475 2.595 5.735 3.195 ;
        RECT  5.370 2.595 5.475 3.025 ;
        RECT  4.750 2.655 5.370 3.025 ;
        RECT  4.655 2.595 4.750 3.025 ;
        RECT  4.395 2.595 4.655 3.195 ;
        RECT  3.575 2.655 4.395 3.025 ;
        RECT  3.315 2.595 3.575 3.195 ;
        RECT  1.085 2.655 3.315 3.025 ;
        RECT  2.815 0.585 3.135 0.895 ;
        RECT  1.705 0.500 2.815 0.895 ;
        END
        ANTENNADIFFAREA     3.9312 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.335 1.885 8.495 2.325 ;
        RECT  5.670 2.165 8.335 2.325 ;
        RECT  5.565 2.110 5.670 2.325 ;
        RECT  5.305 1.885 5.565 2.325 ;
        RECT  2.925 2.165 5.305 2.325 ;
        RECT  2.665 1.885 2.925 2.325 ;
        RECT  2.635 2.110 2.665 2.325 ;
        RECT  2.425 2.110 2.635 2.435 ;
        RECT  0.990 2.275 2.425 2.435 ;
        RECT  0.830 1.510 0.990 2.435 ;
        RECT  0.730 1.510 0.830 1.770 ;
        END
        ANTENNAGATEAREA     1.2922 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.365 1.565 7.465 1.825 ;
        RECT  7.205 1.565 7.365 1.985 ;
        RECT  6.475 1.825 7.205 1.985 ;
        RECT  6.375 1.725 6.475 1.985 ;
        RECT  6.215 1.545 6.375 1.985 ;
        RECT  4.935 1.545 6.215 1.705 ;
        RECT  4.775 1.545 4.935 1.985 ;
        RECT  4.675 1.725 4.775 1.985 ;
        RECT  3.405 1.825 4.675 1.985 ;
        RECT  3.305 1.725 3.405 1.985 ;
        RECT  3.145 1.545 3.305 1.985 ;
        RECT  2.615 1.545 3.145 1.705 ;
        RECT  2.355 1.455 2.615 1.705 ;
        RECT  2.175 1.545 2.355 1.705 ;
        RECT  1.990 1.545 2.175 2.095 ;
        RECT  1.965 1.700 1.990 2.095 ;
        RECT  1.225 1.935 1.965 2.095 ;
        END
        ANTENNAGATEAREA     1.2922 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.815 1.485 6.955 1.645 ;
        RECT  6.655 1.205 6.815 1.645 ;
        RECT  4.290 1.205 6.655 1.365 ;
        RECT  3.990 1.205 4.290 1.615 ;
        RECT  2.955 1.205 3.990 1.365 ;
        RECT  2.795 1.115 2.955 1.365 ;
        RECT  1.745 1.115 2.795 1.275 ;
        RECT  1.505 1.115 1.745 1.665 ;
        END
        ANTENNAGATEAREA     1.2922 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.145 -0.250 9.200 0.250 ;
        RECT  7.885 -0.250 8.145 0.405 ;
        RECT  5.615 -0.250 7.885 0.250 ;
        RECT  5.355 -0.250 5.615 0.405 ;
        RECT  3.295 -0.250 5.355 0.250 ;
        RECT  3.035 -0.250 3.295 0.405 ;
        RECT  0.805 -0.250 3.035 0.250 ;
        RECT  0.545 -0.250 0.805 1.135 ;
        RECT  0.000 -0.250 0.545 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.435 3.440 9.200 3.940 ;
        RECT  8.175 3.285 8.435 3.940 ;
        RECT  7.355 3.440 8.175 3.940 ;
        RECT  7.095 3.285 7.355 3.940 ;
        RECT  6.275 3.440 7.095 3.940 ;
        RECT  6.015 3.285 6.275 3.940 ;
        RECT  5.195 3.440 6.015 3.940 ;
        RECT  4.935 3.285 5.195 3.940 ;
        RECT  4.115 3.440 4.935 3.940 ;
        RECT  3.855 3.285 4.115 3.940 ;
        RECT  3.000 3.440 3.855 3.940 ;
        RECT  2.740 3.285 3.000 3.940 ;
        RECT  1.885 3.440 2.740 3.940 ;
        RECT  1.625 3.285 1.885 3.940 ;
        RECT  0.805 3.440 1.625 3.940 ;
        RECT  0.545 2.875 0.805 3.940 ;
        RECT  0.000 3.440 0.545 3.940 ;
        END
    END VDD
END NAND3X8

MACRO NAND3X6
    CLASS CORE ;
    FOREIGN NAND3X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.675 0.585 6.775 3.155 ;
        RECT  6.415 0.585 6.675 3.195 ;
        RECT  5.005 0.585 6.415 0.885 ;
        RECT  6.105 2.110 6.415 2.810 ;
        RECT  5.670 2.530 6.105 2.790 ;
        RECT  5.515 2.530 5.670 2.810 ;
        RECT  5.255 2.530 5.515 3.195 ;
        RECT  5.185 2.530 5.255 2.995 ;
        RECT  4.495 2.530 5.185 2.790 ;
        RECT  4.745 0.575 5.005 1.175 ;
        RECT  1.905 0.585 4.745 0.885 ;
        RECT  4.235 2.530 4.495 3.195 ;
        RECT  1.085 2.635 4.235 2.935 ;
        END
        ANTENNADIFFAREA     3.5292 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.995 1.405 6.165 1.665 ;
        RECT  5.835 1.405 5.995 1.955 ;
        RECT  5.485 1.795 5.835 1.955 ;
        RECT  5.325 1.795 5.485 2.345 ;
        RECT  3.725 2.185 5.325 2.345 ;
        RECT  3.645 1.810 3.725 2.345 ;
        RECT  3.465 1.810 3.645 2.415 ;
        RECT  3.345 2.110 3.465 2.415 ;
        RECT  1.175 2.255 3.345 2.415 ;
        RECT  1.035 1.950 1.175 2.415 ;
        RECT  1.015 1.510 1.035 2.415 ;
        RECT  0.875 1.510 1.015 2.110 ;
        RECT  0.775 1.510 0.875 1.770 ;
        END
        ANTENNAGATEAREA     0.9360 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.025 1.455 5.655 1.615 ;
        RECT  4.865 1.455 5.025 2.005 ;
        RECT  4.205 1.845 4.865 2.005 ;
        RECT  4.045 1.445 4.205 2.005 ;
        RECT  3.945 1.445 4.045 1.705 ;
        RECT  2.815 1.445 3.945 1.605 ;
        RECT  2.635 1.445 2.815 1.705 ;
        RECT  2.425 1.445 2.635 2.005 ;
        RECT  1.515 1.845 2.425 2.005 ;
        RECT  1.355 1.510 1.515 2.005 ;
        RECT  1.255 1.510 1.355 1.770 ;
        END
        ANTENNAGATEAREA     0.9360 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.555 1.405 4.685 1.665 ;
        RECT  4.395 1.105 4.555 1.665 ;
        RECT  2.175 1.105 4.395 1.265 ;
        RECT  2.015 1.105 2.175 1.580 ;
        RECT  1.995 1.290 2.015 1.580 ;
        RECT  1.735 1.290 1.995 1.665 ;
        END
        ANTENNAGATEAREA     0.9360 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.365 -0.250 6.900 0.250 ;
        RECT  6.105 -0.250 6.365 0.405 ;
        RECT  3.495 -0.250 6.105 0.250 ;
        RECT  3.235 -0.250 3.495 0.405 ;
        RECT  0.835 -0.250 3.235 0.250 ;
        RECT  0.575 -0.250 0.835 1.200 ;
        RECT  0.000 -0.250 0.575 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.115 3.440 6.900 3.940 ;
        RECT  5.855 3.285 6.115 3.940 ;
        RECT  5.005 3.440 5.855 3.940 ;
        RECT  4.745 2.985 5.005 3.940 ;
        RECT  3.900 3.440 4.745 3.940 ;
        RECT  3.280 3.285 3.900 3.940 ;
        RECT  1.955 3.440 3.280 3.940 ;
        RECT  1.695 3.285 1.955 3.940 ;
        RECT  0.805 3.440 1.695 3.940 ;
        RECT  0.545 2.555 0.805 3.940 ;
        RECT  0.000 3.440 0.545 3.940 ;
        END
    END VDD
END NAND3X6

MACRO NAND3X4
    CLASS CORE ;
    FOREIGN NAND3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.290 0.965 4.475 2.465 ;
        RECT  4.235 0.880 4.290 2.465 ;
        RECT  4.210 0.880 4.235 1.205 ;
        RECT  4.015 2.225 4.235 2.465 ;
        RECT  3.950 0.585 4.210 1.205 ;
        RECT  3.935 2.225 4.015 2.585 ;
        RECT  0.875 0.585 3.950 0.825 ;
        RECT  3.675 2.225 3.935 2.960 ;
        RECT  0.875 2.195 2.610 2.455 ;
        RECT  0.635 0.585 0.875 2.455 ;
        RECT  0.585 1.515 0.635 2.175 ;
        END
        ANTENNADIFFAREA     2.7656 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 1.685 3.050 1.945 ;
        RECT  2.790 1.685 2.950 2.795 ;
        RECT  0.335 2.635 2.790 2.795 ;
        RECT  0.335 1.740 0.370 2.000 ;
        RECT  0.160 1.700 0.335 2.795 ;
        RECT  0.125 1.700 0.160 2.585 ;
        RECT  0.110 1.740 0.125 2.180 ;
        END
        ANTENNAGATEAREA     0.5954 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.400 1.795 3.530 2.005 ;
        RECT  3.240 1.345 3.400 2.005 ;
        RECT  2.265 1.345 3.240 1.505 ;
        RECT  2.105 1.345 2.265 2.015 ;
        RECT  1.965 1.700 2.105 2.015 ;
        RECT  1.215 1.855 1.965 2.015 ;
        RECT  1.055 1.745 1.215 2.015 ;
        END
        ANTENNAGATEAREA     0.5954 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.750 1.415 4.010 1.675 ;
        RECT  3.740 1.415 3.750 1.575 ;
        RECT  3.580 1.005 3.740 1.575 ;
        RECT  1.745 1.005 3.580 1.165 ;
        RECT  1.585 1.005 1.745 1.675 ;
        RECT  1.505 1.290 1.585 1.675 ;
        RECT  1.485 1.415 1.505 1.675 ;
        END
        ANTENNAGATEAREA     0.5954 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.905 -0.250 4.600 0.250 ;
        RECT  2.645 -0.250 2.905 0.405 ;
        RECT  0.455 -0.250 2.645 0.250 ;
        RECT  0.195 -0.250 0.455 1.155 ;
        RECT  0.000 -0.250 0.195 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 3.440 4.600 3.940 ;
        RECT  4.215 2.895 4.475 3.940 ;
        RECT  3.395 3.440 4.215 3.940 ;
        RECT  3.135 2.555 3.395 3.940 ;
        RECT  1.465 3.440 3.135 3.940 ;
        RECT  1.205 3.285 1.465 3.940 ;
        RECT  0.385 3.440 1.205 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND3X4

MACRO NAND3X2
    CLASS CORE ;
    FOREIGN NAND3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.110 2.635 2.400 ;
        RECT  0.850 2.135 2.425 2.400 ;
        RECT  1.435 0.475 1.695 1.075 ;
        RECT  0.850 0.915 1.435 1.075 ;
        RECT  0.690 0.915 0.850 2.400 ;
        END
        ANTENNADIFFAREA     1.2729 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.980 1.925 3.095 2.765 ;
        RECT  2.820 1.455 2.980 2.765 ;
        RECT  2.660 1.455 2.820 1.715 ;
        RECT  0.610 2.605 2.820 2.765 ;
        RECT  0.510 2.585 0.610 2.765 ;
        RECT  0.350 1.510 0.510 2.765 ;
        RECT  0.250 1.510 0.350 1.990 ;
        RECT  0.125 1.700 0.250 1.990 ;
        END
        ANTENNAGATEAREA     0.3341 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.245 1.405 2.440 1.665 ;
        RECT  2.085 1.405 2.245 1.955 ;
        RECT  1.295 1.795 2.085 1.955 ;
        RECT  1.255 1.525 1.295 1.955 ;
        RECT  1.045 1.290 1.255 1.955 ;
        RECT  1.035 1.355 1.045 1.955 ;
        END
        ANTENNAGATEAREA     0.3341 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.255 1.875 1.615 ;
        END
        ANTENNAGATEAREA     0.3341 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.090 -0.250 3.220 0.250 ;
        RECT  2.830 -0.250 3.090 1.275 ;
        RECT  0.475 -0.250 2.830 0.250 ;
        RECT  0.215 -0.250 0.475 1.075 ;
        RECT  0.000 -0.250 0.215 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.545 3.440 3.220 3.940 ;
        RECT  1.285 2.945 1.545 3.940 ;
        RECT  0.385 3.440 1.285 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND3X2

MACRO NAND3X1
    CLASS CORE ;
    FOREIGN NAND3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 0.525 1.725 3.135 ;
        RECT  1.435 0.525 1.565 1.125 ;
        RECT  1.505 2.110 1.565 3.135 ;
        RECT  0.785 2.170 1.505 2.330 ;
        RECT  1.435 2.875 1.505 3.135 ;
        RECT  0.525 2.170 0.785 2.430 ;
        END
        ANTENNADIFFAREA     0.9423 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.445 0.375 1.990 ;
        END
        ANTENNAGATEAREA     0.1703 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.480 0.905 1.990 ;
        END
        ANTENNAGATEAREA     0.1703 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.555 1.385 1.815 ;
        RECT  1.250 0.880 1.255 1.170 ;
        RECT  1.090 0.880 1.250 1.815 ;
        RECT  1.045 0.880 1.090 1.170 ;
        END
        ANTENNAGATEAREA     0.1703 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.250 1.840 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 3.440 1.840 3.940 ;
        RECT  0.635 2.895 0.895 3.940 ;
        RECT  0.385 3.440 0.635 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND3X1

MACRO NAND3XL
    CLASS CORE ;
    FOREIGN NAND3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.710 2.110 1.715 3.140 ;
        RECT  1.550 0.820 1.710 3.140 ;
        RECT  1.450 0.820 1.550 1.080 ;
        RECT  1.505 2.110 1.550 3.140 ;
        RECT  1.455 2.235 1.505 3.140 ;
        RECT  0.785 2.235 1.455 2.395 ;
        RECT  0.525 2.235 0.785 2.500 ;
        END
        ANTENNADIFFAREA     0.5824 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.375 0.375 1.990 ;
        END
        ANTENNAGATEAREA     0.0910 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.370 0.835 1.990 ;
        END
        ANTENNAGATEAREA     0.0910 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.345 1.350 1.890 ;
        RECT  1.045 1.345 1.255 1.990 ;
        END
        ANTENNAGATEAREA     0.0910 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.250 1.840 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 3.440 1.840 3.940 ;
        RECT  0.635 2.890 0.895 3.940 ;
        RECT  0.385 3.440 0.635 3.940 ;
        RECT  0.125 2.890 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND3XL

MACRO NAND2X8
    CLASS CORE ;
    FOREIGN NAND2X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.125 1.700 5.395 2.590 ;
        RECT  4.750 0.900 5.125 2.590 ;
        RECT  4.725 0.880 4.750 2.590 ;
        RECT  4.605 0.880 4.725 1.300 ;
        RECT  4.015 2.190 4.725 2.590 ;
        RECT  4.275 0.585 4.605 1.300 ;
        RECT  0.945 0.585 4.275 0.985 ;
        RECT  3.955 2.190 4.015 2.995 ;
        RECT  3.695 2.190 3.955 3.140 ;
        RECT  2.935 2.190 3.695 2.590 ;
        RECT  2.675 2.190 2.935 3.140 ;
        RECT  1.915 2.190 2.675 2.590 ;
        RECT  1.655 2.190 1.915 3.140 ;
        RECT  0.895 2.190 1.655 2.590 ;
        RECT  0.635 2.190 0.895 3.140 ;
        RECT  0.585 2.745 0.635 2.995 ;
        END
        ANTENNADIFFAREA     2.7480 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.295 1.315 3.555 1.615 ;
        RECT  2.055 1.315 3.295 1.475 ;
        RECT  1.690 1.315 2.055 1.615 ;
        RECT  0.555 1.315 1.690 1.475 ;
        RECT  0.395 1.315 0.555 1.925 ;
        RECT  0.335 1.665 0.395 1.925 ;
        RECT  0.295 1.665 0.335 1.990 ;
        RECT  0.125 1.700 0.295 1.990 ;
        END
        ANTENNAGATEAREA     1.1700 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 1.665 4.435 1.955 ;
        RECT  2.910 1.795 3.990 1.955 ;
        RECT  2.475 1.665 2.910 1.955 ;
        RECT  1.255 1.795 2.475 1.955 ;
        RECT  1.045 1.700 1.255 1.990 ;
        RECT  1.035 1.700 1.045 1.955 ;
        RECT  0.775 1.665 1.035 1.955 ;
        END
        ANTENNAGATEAREA     1.1700 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.755 -0.250 5.520 0.250 ;
        RECT  3.495 -0.250 3.755 0.405 ;
        RECT  2.055 -0.250 3.495 0.250 ;
        RECT  1.795 -0.250 2.055 0.405 ;
        RECT  0.385 -0.250 1.795 0.250 ;
        RECT  0.125 -0.250 0.385 1.095 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 3.440 5.520 3.940 ;
        RECT  4.205 2.935 4.465 3.940 ;
        RECT  3.445 3.440 4.205 3.940 ;
        RECT  3.185 2.895 3.445 3.940 ;
        RECT  2.425 3.440 3.185 3.940 ;
        RECT  2.165 2.935 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.935 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.255 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND2X8

MACRO NAND2X6
    CLASS CORE ;
    FOREIGN NAND2X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.735 0.755 4.035 2.810 ;
        RECT  2.905 0.755 3.735 1.055 ;
        RECT  2.935 2.110 3.735 2.810 ;
        RECT  2.885 2.110 2.935 3.195 ;
        RECT  2.645 0.495 2.905 1.095 ;
        RECT  2.675 2.255 2.885 3.195 ;
        RECT  1.915 2.255 2.675 2.555 ;
        RECT  1.230 0.755 2.645 1.055 ;
        RECT  1.655 2.255 1.915 3.195 ;
        RECT  0.895 2.255 1.655 2.555 ;
        RECT  1.205 0.695 1.230 1.055 ;
        RECT  0.945 0.495 1.205 1.095 ;
        RECT  0.635 2.255 0.895 3.195 ;
        RECT  0.585 2.745 0.635 2.995 ;
        END
        ANTENNADIFFAREA     2.0862 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 1.405 3.555 1.665 ;
        RECT  3.295 1.305 3.460 1.665 ;
        RECT  2.255 1.305 3.295 1.465 ;
        RECT  1.995 1.305 2.255 1.665 ;
        RECT  0.405 1.305 1.995 1.465 ;
        RECT  0.335 1.305 0.405 1.925 ;
        RECT  0.245 1.305 0.335 1.990 ;
        RECT  0.125 1.510 0.245 1.990 ;
        END
        ANTENNAGATEAREA     0.9321 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.645 2.735 1.805 ;
        RECT  2.475 1.645 2.635 2.035 ;
        RECT  1.255 1.875 2.475 2.035 ;
        RECT  0.975 1.645 1.255 2.035 ;
        END
        ANTENNAGATEAREA     0.9321 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.755 -0.250 4.600 0.250 ;
        RECT  3.495 -0.250 3.755 0.405 ;
        RECT  2.055 -0.250 3.495 0.250 ;
        RECT  1.795 -0.250 2.055 0.405 ;
        RECT  0.385 -0.250 1.795 0.250 ;
        RECT  0.125 -0.250 0.385 1.095 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.475 3.440 4.600 3.940 ;
        RECT  3.215 3.285 3.475 3.940 ;
        RECT  2.425 3.440 3.215 3.940 ;
        RECT  2.165 2.895 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.895 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.255 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND2X6

MACRO NAND2X4
    CLASS CORE ;
    FOREIGN NAND2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 0.585 3.110 2.715 ;
        RECT  2.885 0.585 2.910 1.580 ;
        RECT  2.005 2.515 2.910 2.715 ;
        RECT  2.835 0.585 2.885 1.185 ;
        RECT  1.530 0.975 2.835 1.175 ;
        RECT  1.745 2.515 2.005 3.195 ;
        RECT  0.925 2.515 1.745 2.715 ;
        RECT  1.125 0.915 1.530 1.175 ;
        RECT  0.665 2.255 0.925 3.195 ;
        RECT  0.585 2.745 0.665 2.995 ;
        END
        ANTENNADIFFAREA     1.4224 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 1.645 2.145 1.905 ;
        RECT  1.885 1.355 2.045 1.905 ;
        RECT  0.795 1.355 1.885 1.515 ;
        RECT  0.585 1.290 0.795 1.905 ;
        RECT  0.475 1.515 0.585 1.905 ;
        END
        ANTENNAGATEAREA     0.5850 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.700 2.725 2.075 ;
        RECT  2.425 1.700 2.585 2.335 ;
        RECT  1.375 2.175 2.425 2.335 ;
        RECT  1.215 1.715 1.375 2.335 ;
        RECT  1.115 1.715 1.215 1.875 ;
        END
        ANTENNAGATEAREA     0.5850 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.275 -0.250 3.220 0.250 ;
        RECT  2.015 -0.250 2.275 0.795 ;
        RECT  0.535 -0.250 2.015 0.250 ;
        RECT  0.275 -0.250 0.535 1.085 ;
        RECT  0.000 -0.250 0.275 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 3.440 3.220 3.940 ;
        RECT  2.310 2.895 2.570 3.940 ;
        RECT  1.465 3.440 2.310 3.940 ;
        RECT  1.205 2.895 1.465 3.940 ;
        RECT  0.385 3.440 1.205 3.940 ;
        RECT  0.125 2.215 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND2X4

MACRO NAND2X2
    CLASS CORE ;
    FOREIGN NAND2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 1.925 2.175 2.400 ;
        RECT  1.965 1.380 2.125 2.400 ;
        RECT  1.640 1.380 1.965 1.540 ;
        RECT  0.925 2.195 1.965 2.355 ;
        RECT  1.480 0.950 1.640 1.540 ;
        RECT  1.265 0.950 1.480 1.110 ;
        RECT  1.005 0.850 1.265 1.110 ;
        RECT  0.665 2.195 0.925 3.135 ;
        RECT  0.585 2.745 0.665 2.995 ;
        END
        ANTENNADIFFAREA     0.7561 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 1.725 1.785 2.015 ;
        RECT  0.510 1.855 1.575 2.015 ;
        RECT  0.250 1.585 0.510 2.015 ;
        RECT  0.125 1.700 0.250 2.015 ;
        END
        ANTENNAGATEAREA     0.3172 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.065 1.290 1.255 1.580 ;
        RECT  0.805 1.290 1.065 1.675 ;
        END
        ANTENNAGATEAREA     0.3172 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 -0.250 2.300 0.250 ;
        RECT  1.915 -0.250 2.175 1.140 ;
        RECT  0.385 -0.250 1.915 0.250 ;
        RECT  0.125 -0.250 0.385 1.140 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 3.440 2.300 3.940 ;
        RECT  1.205 2.555 1.465 3.940 ;
        RECT  0.385 3.440 1.205 3.940 ;
        RECT  0.125 2.555 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND2X2

MACRO NAND2X1
    CLASS CORE ;
    FOREIGN NAND2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.380 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.035 1.265 2.585 ;
        RECT  1.105 1.035 1.255 2.810 ;
        RECT  0.995 1.035 1.105 1.355 ;
        RECT  1.045 2.275 1.105 2.810 ;
        RECT  0.525 2.275 1.045 2.535 ;
        END
        ANTENNADIFFAREA     0.4404 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.405 1.770 ;
        END
        ANTENNAGATEAREA     0.1586 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.725 0.925 1.985 ;
        RECT  0.635 1.290 0.795 1.985 ;
        RECT  0.585 1.290 0.635 1.765 ;
        END
        ANTENNAGATEAREA     0.1586 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 -0.250 1.380 0.250 ;
        RECT  0.145 -0.250 0.405 1.085 ;
        RECT  0.000 -0.250 0.145 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 3.440 1.380 3.940 ;
        RECT  0.995 3.285 1.255 3.940 ;
        RECT  0.385 3.440 0.995 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND2X1

MACRO NAND2XL
    CLASS CORE ;
    FOREIGN NAND2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.380 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 0.810 1.265 2.455 ;
        RECT  1.045 0.810 1.105 1.170 ;
        RECT  0.785 2.295 1.105 2.455 ;
        RECT  0.995 0.810 1.045 1.070 ;
        RECT  0.525 2.295 0.785 2.555 ;
        END
        ANTENNADIFFAREA     0.2346 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.405 1.770 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.510 0.925 1.990 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.250 1.380 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 3.440 1.380 3.940 ;
        RECT  0.995 2.895 1.255 3.940 ;
        RECT  0.385 3.440 0.995 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END NAND2XL

MACRO MXI3X4
    CLASS CORE ;
    FOREIGN MXI3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.105 1.290 8.155 2.585 ;
        RECT  7.865 0.600 8.105 3.050 ;
        RECT  7.815 0.600 7.865 1.200 ;
        RECT  7.845 2.110 7.865 3.050 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.265 1.925 6.315 2.400 ;
        RECT  6.105 1.490 6.265 2.400 ;
        RECT  5.965 1.490 6.105 1.750 ;
        END
        ANTENNAGATEAREA     0.3731 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.435 2.685 1.695 ;
        RECT  2.425 1.435 2.635 1.990 ;
        END
        ANTENNAGATEAREA     0.2938 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.570 1.950 3.580 2.210 ;
        RECT  3.310 1.700 3.570 2.210 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.260 2.190 1.820 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.535 0.385 2.090 ;
        END
        ANTENNAGATEAREA     0.2158 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.585 -0.250 8.740 0.250 ;
        RECT  8.325 -0.250 8.585 1.095 ;
        RECT  7.520 -0.250 8.325 0.250 ;
        RECT  7.260 -0.250 7.520 0.405 ;
        RECT  6.435 -0.250 7.260 0.250 ;
        RECT  6.175 -0.250 6.435 0.405 ;
        RECT  3.740 -0.250 6.175 0.250 ;
        RECT  3.580 -0.250 3.740 1.130 ;
        RECT  2.505 -0.250 3.580 0.250 ;
        RECT  2.245 -0.250 2.505 1.045 ;
        RECT  0.360 -0.250 2.245 0.250 ;
        RECT  0.200 -0.250 0.360 1.295 ;
        RECT  0.000 -0.250 0.200 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.615 3.440 8.740 3.940 ;
        RECT  8.355 2.205 8.615 3.940 ;
        RECT  7.545 3.440 8.355 3.940 ;
        RECT  7.385 2.200 7.545 3.940 ;
        RECT  6.365 3.440 7.385 3.940 ;
        RECT  6.105 3.285 6.365 3.940 ;
        RECT  3.900 3.440 6.105 3.940 ;
        RECT  3.640 3.285 3.900 3.940 ;
        RECT  2.495 3.440 3.640 3.940 ;
        RECT  2.235 3.090 2.495 3.940 ;
        RECT  0.385 3.440 2.235 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.555 1.470 7.660 1.730 ;
        RECT  7.395 0.615 7.555 1.730 ;
        RECT  4.860 0.615 7.395 0.775 ;
        RECT  7.045 1.535 7.205 3.105 ;
        RECT  6.855 1.535 7.045 1.795 ;
        RECT  5.865 2.945 7.045 3.105 ;
        RECT  6.720 1.000 6.980 1.260 ;
        RECT  6.675 2.070 6.865 2.760 ;
        RECT  6.675 1.100 6.720 1.260 ;
        RECT  6.515 1.100 6.675 2.760 ;
        RECT  5.470 2.600 6.515 2.760 ;
        RECT  5.785 1.025 5.885 1.285 ;
        RECT  5.785 2.090 5.870 2.350 ;
        RECT  5.705 2.945 5.865 3.200 ;
        RECT  5.625 1.025 5.785 2.350 ;
        RECT  4.480 3.040 5.705 3.200 ;
        RECT  5.480 1.395 5.625 1.665 ;
        RECT  5.610 2.090 5.625 2.350 ;
        RECT  5.300 2.600 5.470 2.860 ;
        RECT  5.300 0.955 5.320 1.215 ;
        RECT  5.140 0.955 5.300 2.860 ;
        RECT  5.060 0.955 5.140 1.215 ;
        RECT  4.860 2.110 4.960 2.710 ;
        RECT  4.700 0.615 4.860 2.710 ;
        RECT  4.550 0.695 4.700 1.295 ;
        RECT  4.320 2.940 4.480 3.200 ;
        RECT  4.350 2.090 4.450 2.690 ;
        RECT  4.190 0.575 4.350 2.690 ;
        RECT  2.865 2.940 4.320 3.100 ;
        RECT  4.040 0.575 4.190 1.175 ;
        RECT  3.850 1.360 4.010 2.750 ;
        RECT  3.750 1.360 3.850 1.720 ;
        RECT  3.090 2.590 3.850 2.750 ;
        RECT  3.380 1.360 3.750 1.520 ;
        RECT  3.220 0.515 3.380 1.520 ;
        RECT  2.980 0.515 3.220 0.775 ;
        RECT  2.865 1.035 3.025 2.345 ;
        RECT  2.835 1.955 2.865 2.345 ;
        RECT  2.705 2.710 2.865 3.100 ;
        RECT  2.470 2.185 2.835 2.345 ;
        RECT  1.340 2.710 2.705 2.870 ;
        RECT  2.310 2.185 2.470 2.530 ;
        RECT  1.430 2.370 2.310 2.530 ;
        RECT  1.770 0.780 1.995 1.040 ;
        RECT  1.770 2.030 1.920 2.190 ;
        RECT  1.610 0.780 1.770 2.190 ;
        RECT  1.270 1.605 1.430 2.530 ;
        RECT  1.240 0.695 1.400 1.410 ;
        RECT  1.080 2.710 1.340 2.970 ;
        RECT  1.075 1.250 1.240 1.410 ;
        RECT  1.075 2.710 1.080 2.870 ;
        RECT  0.915 1.250 1.075 2.870 ;
        RECT  0.735 0.790 0.925 1.050 ;
        RECT  0.575 0.790 0.735 2.855 ;
    END
END MXI3X4

MACRO MXI3X2
    CLASS CORE ;
    FOREIGN MXI3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 0.600 7.695 3.050 ;
        RECT  7.435 0.600 7.485 1.200 ;
        RECT  7.435 2.110 7.485 3.050 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.265 1.290 6.315 1.580 ;
        RECT  6.105 1.290 6.265 1.680 ;
        RECT  6.015 1.520 6.105 1.680 ;
        RECT  5.755 1.520 6.015 1.780 ;
        END
        ANTENNAGATEAREA     0.2951 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.435 2.685 1.695 ;
        RECT  2.425 1.435 2.635 1.990 ;
        END
        ANTENNAGATEAREA     0.2275 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.465 1.700 3.555 1.990 ;
        RECT  3.205 1.700 3.465 2.210 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 1.250 2.235 1.635 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.600 0.385 2.155 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.145 -0.250 7.820 0.250 ;
        RECT  6.885 -0.250 7.145 0.405 ;
        RECT  6.225 -0.250 6.885 0.250 ;
        RECT  5.965 -0.250 6.225 0.405 ;
        RECT  3.715 -0.250 5.965 0.250 ;
        RECT  3.455 -0.250 3.715 0.405 ;
        RECT  2.370 -0.250 3.455 0.250 ;
        RECT  2.110 -0.250 2.370 1.035 ;
        RECT  0.385 -0.250 2.110 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.145 3.440 7.820 3.940 ;
        RECT  6.885 2.850 7.145 3.940 ;
        RECT  6.160 3.440 6.885 3.940 ;
        RECT  5.900 3.285 6.160 3.940 ;
        RECT  3.675 3.440 5.900 3.940 ;
        RECT  3.415 3.285 3.675 3.940 ;
        RECT  2.445 3.440 3.415 3.940 ;
        RECT  2.285 2.985 2.445 3.940 ;
        RECT  0.385 3.440 2.285 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.120 1.470 7.260 1.730 ;
        RECT  6.960 0.625 7.120 1.730 ;
        RECT  5.705 0.625 6.960 0.785 ;
        RECT  6.660 1.000 6.775 1.260 ;
        RECT  6.660 1.955 6.710 2.555 ;
        RECT  6.610 1.000 6.660 2.555 ;
        RECT  6.365 2.945 6.630 3.215 ;
        RECT  6.500 1.000 6.610 2.685 ;
        RECT  6.450 1.955 6.500 2.685 ;
        RECT  5.265 2.525 6.450 2.685 ;
        RECT  5.605 2.945 6.365 3.105 ;
        RECT  5.745 1.035 5.795 1.295 ;
        RECT  5.575 1.030 5.745 1.295 ;
        RECT  5.545 0.540 5.705 0.785 ;
        RECT  5.575 2.085 5.670 2.345 ;
        RECT  5.445 2.945 5.605 3.260 ;
        RECT  5.415 1.030 5.575 2.345 ;
        RECT  4.775 0.540 5.545 0.700 ;
        RECT  4.770 3.100 5.445 3.260 ;
        RECT  5.410 1.405 5.415 2.345 ;
        RECT  5.305 1.405 5.410 1.665 ;
        RECT  5.120 2.525 5.265 2.885 ;
        RECT  5.120 0.965 5.235 1.225 ;
        RECT  4.960 0.965 5.120 2.885 ;
        RECT  4.705 0.540 4.775 1.290 ;
        RECT  4.610 2.945 4.770 3.260 ;
        RECT  4.705 2.425 4.755 2.685 ;
        RECT  4.545 0.540 4.705 2.685 ;
        RECT  2.795 2.945 4.610 3.105 ;
        RECT  4.515 0.540 4.545 1.290 ;
        RECT  4.495 2.425 4.545 2.685 ;
        RECT  4.145 0.850 4.305 2.765 ;
        RECT  4.005 0.850 4.145 1.110 ;
        RECT  3.985 2.510 4.145 2.765 ;
        RECT  3.805 1.360 3.940 2.330 ;
        RECT  3.780 1.360 3.805 2.740 ;
        RECT  3.770 1.360 3.780 1.520 ;
        RECT  3.645 2.170 3.780 2.740 ;
        RECT  3.610 0.625 3.770 1.520 ;
        RECT  2.980 2.580 3.645 2.740 ;
        RECT  3.135 0.625 3.610 0.785 ;
        RECT  2.875 0.445 3.135 0.785 ;
        RECT  2.865 0.975 3.025 2.385 ;
        RECT  2.680 0.975 2.865 1.235 ;
        RECT  2.835 2.015 2.865 2.385 ;
        RECT  2.240 2.225 2.835 2.385 ;
        RECT  2.635 2.630 2.795 3.105 ;
        RECT  1.340 2.630 2.635 2.790 ;
        RECT  2.080 1.925 2.240 2.385 ;
        RECT  1.755 1.925 2.080 2.085 ;
        RECT  1.415 2.270 1.895 2.430 ;
        RECT  1.705 0.780 1.860 1.040 ;
        RECT  1.595 1.815 1.755 2.085 ;
        RECT  1.545 0.780 1.705 1.585 ;
        RECT  1.415 1.425 1.545 1.585 ;
        RECT  1.255 1.425 1.415 2.430 ;
        RECT  1.090 0.880 1.350 1.140 ;
        RECT  1.080 2.630 1.340 2.890 ;
        RECT  1.075 0.980 1.090 1.140 ;
        RECT  1.075 2.630 1.080 2.790 ;
        RECT  0.915 0.980 1.075 2.790 ;
        RECT  0.575 0.870 0.735 2.855 ;
    END
END MXI3X2

MACRO MXI3X1
    CLASS CORE ;
    FOREIGN MXI3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.080 0.520 7.240 3.025 ;
        RECT  7.020 0.520 7.080 0.780 ;
        RECT  7.025 2.335 7.080 3.025 ;
        RECT  6.975 2.765 7.025 3.025 ;
        END
        ANTENNADIFFAREA     0.3264 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.755 6.860 1.985 ;
        RECT  6.565 1.700 6.775 1.990 ;
        RECT  6.310 1.755 6.565 1.985 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 2.880 0.935 3.240 ;
        END
        ANTENNAGATEAREA     0.1313 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.200 1.695 3.555 2.090 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.290 2.635 1.610 ;
        RECT  2.290 1.380 2.425 1.610 ;
        RECT  2.030 1.380 2.290 1.660 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.635 0.390 1.895 ;
        RECT  0.130 1.290 0.335 1.895 ;
        RECT  0.125 1.290 0.130 1.765 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.680 -0.250 7.360 0.250 ;
        RECT  6.420 -0.250 6.680 0.405 ;
        RECT  5.820 -0.250 6.420 0.250 ;
        RECT  5.660 -0.250 5.820 0.815 ;
        RECT  3.620 -0.250 5.660 0.250 ;
        RECT  3.360 -0.250 3.620 0.405 ;
        RECT  2.465 -0.250 3.360 0.250 ;
        RECT  2.205 -0.250 2.465 1.090 ;
        RECT  0.385 -0.250 2.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 3.440 7.360 3.940 ;
        RECT  6.465 2.805 6.725 3.940 ;
        RECT  6.095 3.440 6.465 3.940 ;
        RECT  5.935 2.700 6.095 3.940 ;
        RECT  3.830 3.440 5.935 3.940 ;
        RECT  3.570 3.285 3.830 3.940 ;
        RECT  2.365 3.440 3.570 3.940 ;
        RECT  2.105 3.105 2.365 3.940 ;
        RECT  0.385 3.440 2.105 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.840 1.100 6.900 1.360 ;
        RECT  6.680 0.730 6.840 1.360 ;
        RECT  6.160 0.730 6.680 0.890 ;
        RECT  6.095 2.170 6.680 2.330 ;
        RECT  6.340 1.085 6.500 1.525 ;
        RECT  6.095 1.345 6.340 1.525 ;
        RECT  6.000 0.730 6.160 1.160 ;
        RECT  5.935 1.345 6.095 2.330 ;
        RECT  5.480 1.000 6.000 1.160 ;
        RECT  5.210 1.585 5.935 1.845 ;
        RECT  5.565 2.070 5.725 3.105 ;
        RECT  2.810 2.945 5.565 3.105 ;
        RECT  5.320 0.510 5.480 1.160 ;
        RECT  5.225 2.040 5.385 2.700 ;
        RECT  4.675 0.510 5.320 0.670 ;
        RECT  5.030 2.040 5.225 2.200 ;
        RECT  5.030 0.850 5.135 1.110 ;
        RECT  4.870 0.850 5.030 2.200 ;
        RECT  4.675 2.420 4.925 2.680 ;
        RECT  4.515 0.510 4.675 2.680 ;
        RECT  4.415 0.830 4.515 1.090 ;
        RECT  4.235 2.280 4.320 2.540 ;
        RECT  4.075 0.845 4.235 2.540 ;
        RECT  3.905 0.845 4.075 1.105 ;
        RECT  3.735 1.320 3.895 2.440 ;
        RECT  3.480 1.320 3.735 1.480 ;
        RECT  3.340 2.280 3.735 2.440 ;
        RECT  3.320 0.615 3.480 1.480 ;
        RECT  3.080 2.280 3.340 2.540 ;
        RECT  3.040 0.615 3.320 0.775 ;
        RECT  2.780 0.515 3.040 0.775 ;
        RECT  2.830 1.030 2.990 2.010 ;
        RECT  2.570 1.850 2.830 2.570 ;
        RECT  2.650 2.760 2.810 3.105 ;
        RECT  1.400 2.760 2.650 2.920 ;
        RECT  1.760 1.850 2.570 2.010 ;
        RECT  1.675 1.030 1.835 1.480 ;
        RECT  1.695 2.420 1.795 2.580 ;
        RECT  1.600 1.720 1.760 2.010 ;
        RECT  1.535 2.190 1.695 2.580 ;
        RECT  1.415 1.320 1.675 1.480 ;
        RECT  1.415 2.190 1.535 2.350 ;
        RECT  1.365 0.455 1.465 0.715 ;
        RECT  1.255 1.320 1.415 2.350 ;
        RECT  1.280 2.760 1.400 3.240 ;
        RECT  1.205 0.455 1.365 1.140 ;
        RECT  1.120 2.540 1.280 3.240 ;
        RECT  1.075 0.980 1.205 1.140 ;
        RECT  1.075 2.540 1.120 2.700 ;
        RECT  0.915 0.980 1.075 2.700 ;
        RECT  0.735 0.500 0.905 0.760 ;
        RECT  0.575 0.500 0.735 2.580 ;
    END
END MXI3X1

MACRO MXI3XL
    CLASS CORE ;
    FOREIGN MXI3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 0.510 7.240 2.680 ;
        RECT  7.080 0.510 7.235 2.935 ;
        RECT  7.050 0.510 7.080 0.945 ;
        RECT  7.025 2.335 7.080 2.935 ;
        RECT  7.025 0.510 7.050 0.770 ;
        RECT  6.975 2.675 7.025 2.935 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.755 6.860 1.985 ;
        RECT  6.565 1.700 6.775 1.990 ;
        RECT  6.310 1.755 6.565 1.985 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 2.880 0.960 3.220 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.200 1.700 3.555 2.090 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.290 2.635 1.615 ;
        RECT  2.315 1.385 2.425 1.615 ;
        RECT  2.055 1.385 2.315 1.665 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.635 0.390 1.895 ;
        RECT  0.130 1.290 0.335 1.895 ;
        RECT  0.125 1.290 0.130 1.765 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.655 -0.250 7.360 0.250 ;
        RECT  6.395 -0.250 6.655 0.405 ;
        RECT  5.815 -0.250 6.395 0.250 ;
        RECT  5.655 -0.250 5.815 0.815 ;
        RECT  3.620 -0.250 5.655 0.250 ;
        RECT  3.360 -0.250 3.620 0.405 ;
        RECT  2.465 -0.250 3.360 0.250 ;
        RECT  2.205 -0.250 2.465 1.095 ;
        RECT  0.385 -0.250 2.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.800 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 3.440 7.360 3.940 ;
        RECT  6.465 2.655 6.725 3.940 ;
        RECT  6.070 3.440 6.465 3.940 ;
        RECT  5.910 2.700 6.070 3.940 ;
        RECT  3.830 3.440 5.910 3.940 ;
        RECT  3.570 3.285 3.830 3.940 ;
        RECT  2.385 3.440 3.570 3.940 ;
        RECT  2.125 3.105 2.385 3.940 ;
        RECT  0.385 3.440 2.125 3.940 ;
        RECT  0.125 2.860 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.835 1.020 6.870 1.280 ;
        RECT  6.675 0.630 6.835 1.280 ;
        RECT  6.095 2.170 6.680 2.330 ;
        RECT  6.155 0.630 6.675 0.790 ;
        RECT  6.335 0.970 6.495 1.525 ;
        RECT  6.095 1.345 6.335 1.525 ;
        RECT  5.995 0.630 6.155 1.160 ;
        RECT  5.935 1.345 6.095 2.330 ;
        RECT  5.475 1.000 5.995 1.160 ;
        RECT  5.210 1.605 5.935 1.865 ;
        RECT  5.730 2.090 5.755 2.350 ;
        RECT  5.570 2.090 5.730 3.050 ;
        RECT  3.705 2.890 5.570 3.050 ;
        RECT  5.315 0.480 5.475 1.160 ;
        RECT  5.225 2.075 5.385 2.700 ;
        RECT  4.660 0.480 5.315 0.640 ;
        RECT  5.005 2.075 5.225 2.235 ;
        RECT  5.005 0.820 5.135 1.425 ;
        RECT  4.975 0.820 5.005 2.235 ;
        RECT  4.845 1.265 4.975 2.235 ;
        RECT  4.665 2.415 4.925 2.675 ;
        RECT  4.660 2.415 4.665 2.575 ;
        RECT  4.500 0.480 4.660 2.575 ;
        RECT  4.465 0.820 4.500 1.080 ;
        RECT  4.245 2.415 4.320 2.675 ;
        RECT  4.165 0.920 4.245 2.675 ;
        RECT  4.085 0.820 4.165 2.675 ;
        RECT  3.905 0.820 4.085 1.080 ;
        RECT  3.745 1.260 3.905 2.455 ;
        RECT  3.630 1.260 3.745 1.520 ;
        RECT  3.340 2.295 3.745 2.455 ;
        RECT  3.545 2.765 3.705 3.050 ;
        RECT  3.480 1.260 3.630 1.420 ;
        RECT  1.405 2.765 3.545 2.925 ;
        RECT  3.320 0.615 3.480 1.420 ;
        RECT  3.080 2.295 3.340 2.555 ;
        RECT  3.040 0.615 3.320 0.775 ;
        RECT  2.780 0.515 3.040 0.775 ;
        RECT  2.830 1.035 2.990 2.005 ;
        RECT  2.570 1.845 2.830 2.570 ;
        RECT  1.785 1.845 2.570 2.005 ;
        RECT  1.755 1.035 1.855 1.295 ;
        RECT  1.545 2.185 1.805 2.525 ;
        RECT  1.625 1.745 1.785 2.005 ;
        RECT  1.595 1.035 1.755 1.480 ;
        RECT  1.445 1.320 1.595 1.480 ;
        RECT  1.445 2.185 1.545 2.345 ;
        RECT  1.365 0.455 1.465 0.715 ;
        RECT  1.285 1.320 1.445 2.345 ;
        RECT  1.300 2.765 1.405 3.215 ;
        RECT  1.205 0.455 1.365 1.140 ;
        RECT  1.140 2.525 1.300 3.215 ;
        RECT  1.105 0.980 1.205 1.140 ;
        RECT  1.105 2.525 1.140 2.685 ;
        RECT  0.945 0.980 1.105 2.685 ;
        RECT  0.765 0.455 0.905 0.715 ;
        RECT  0.605 0.455 0.765 2.525 ;
    END
END MXI3XL

MACRO MX3X4
    CLASS CORE ;
    FOREIGN MX3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.280 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.760 1.285 8.155 1.995 ;
        RECT  7.695 0.595 7.760 2.585 ;
        RECT  7.645 0.595 7.695 2.995 ;
        RECT  7.520 0.595 7.645 3.105 ;
        RECT  7.385 0.595 7.520 0.855 ;
        RECT  7.385 2.165 7.520 3.105 ;
        END
        ANTENNADIFFAREA     0.8026 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.765 2.110 6.775 2.400 ;
        RECT  6.505 1.855 6.765 2.400 ;
        RECT  6.305 2.240 6.505 2.400 ;
        RECT  6.145 2.240 6.305 2.745 ;
        RECT  4.685 2.585 6.145 2.745 ;
        END
        ANTENNAGATEAREA     0.3848 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 2.540 3.255 2.800 ;
        RECT  2.885 2.520 3.095 2.810 ;
        RECT  1.135 2.575 2.885 2.735 ;
        RECT  2.370 0.505 2.630 0.765 ;
        RECT  1.040 0.605 2.370 0.765 ;
        RECT  1.135 1.480 1.210 1.740 ;
        RECT  1.040 1.480 1.135 2.735 ;
        RECT  0.975 0.605 1.040 2.735 ;
        RECT  0.880 0.605 0.975 1.740 ;
        END
        ANTENNAGATEAREA     0.3861 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 2.110 0.795 2.400 ;
        RECT  0.540 1.575 0.700 2.400 ;
        RECT  0.505 1.575 0.540 1.835 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.780 1.290 2.240 1.625 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.290 4.475 1.810 ;
        RECT  4.060 1.550 4.265 1.810 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.105 -0.250 8.280 0.250 ;
        RECT  7.945 -0.250 8.105 1.075 ;
        RECT  7.135 -0.250 7.945 0.250 ;
        RECT  6.875 -0.250 7.135 0.805 ;
        RECT  4.470 -0.250 6.875 0.250 ;
        RECT  4.210 -0.250 4.470 0.405 ;
        RECT  1.820 -0.250 4.210 0.250 ;
        RECT  1.560 -0.250 1.820 0.405 ;
        RECT  1.010 -0.250 1.560 0.340 ;
        RECT  0.750 -0.250 1.010 0.415 ;
        RECT  0.000 -0.250 0.750 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.105 3.440 8.280 3.940 ;
        RECT  7.945 2.275 8.105 3.940 ;
        RECT  7.135 3.440 7.945 3.940 ;
        RECT  6.875 2.955 7.135 3.940 ;
        RECT  4.565 3.440 6.875 3.940 ;
        RECT  4.305 3.285 4.565 3.940 ;
        RECT  1.925 3.440 4.305 3.940 ;
        RECT  1.665 3.285 1.925 3.940 ;
        RECT  0.980 3.355 1.665 3.940 ;
        RECT  0.720 3.275 0.980 3.940 ;
        RECT  0.000 3.440 0.720 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.175 1.035 7.335 1.980 ;
        RECT  6.625 1.035 7.175 1.195 ;
        RECT  7.015 1.820 7.175 2.770 ;
        RECT  6.650 2.610 7.015 2.770 ;
        RECT  6.830 1.375 6.990 1.635 ;
        RECT  6.115 1.475 6.830 1.635 ;
        RECT  6.500 2.610 6.650 3.155 ;
        RECT  6.365 0.580 6.625 1.195 ;
        RECT  6.490 2.610 6.500 3.205 ;
        RECT  6.240 2.945 6.490 3.205 ;
        RECT  3.865 2.945 6.240 3.105 ;
        RECT  5.940 0.675 6.115 1.635 ;
        RECT  5.855 0.675 5.940 2.360 ;
        RECT  5.780 1.475 5.855 2.360 ;
        RECT  5.555 0.535 5.605 1.135 ;
        RECT  5.395 0.535 5.555 2.320 ;
        RECT  5.345 0.535 5.395 1.135 ;
        RECT  5.220 2.060 5.395 2.320 ;
        RECT  3.400 0.590 5.345 0.750 ;
        RECT  5.020 1.265 5.210 1.525 ;
        RECT  4.970 0.930 5.020 1.525 ;
        RECT  4.810 0.930 4.970 2.215 ;
        RECT  4.760 0.930 4.810 1.090 ;
        RECT  4.710 1.955 4.810 2.215 ;
        RECT  3.835 2.075 4.025 2.675 ;
        RECT  3.835 0.975 3.910 1.235 ;
        RECT  3.705 2.945 3.865 3.220 ;
        RECT  3.765 0.975 3.835 2.675 ;
        RECT  3.675 0.975 3.765 2.455 ;
        RECT  2.345 3.060 3.705 3.220 ;
        RECT  3.650 0.975 3.675 1.235 ;
        RECT  3.365 2.050 3.465 2.310 ;
        RECT  3.365 0.590 3.400 1.190 ;
        RECT  3.205 0.590 3.365 2.310 ;
        RECT  3.140 0.590 3.205 1.190 ;
        RECT  2.800 0.945 2.960 2.340 ;
        RECT  2.175 0.945 2.800 1.105 ;
        RECT  2.225 2.180 2.800 2.340 ;
        RECT  2.460 1.540 2.620 1.995 ;
        RECT  1.560 1.825 2.460 1.995 ;
        RECT  2.185 2.935 2.345 3.220 ;
        RECT  0.335 2.935 2.185 3.095 ;
        RECT  1.400 1.135 1.560 2.250 ;
        RECT  1.380 1.135 1.400 1.295 ;
        RECT  1.320 1.990 1.400 2.250 ;
        RECT  1.220 1.035 1.380 1.295 ;
        RECT  0.310 0.600 0.445 1.200 ;
        RECT  0.310 2.155 0.335 3.095 ;
        RECT  0.185 0.600 0.310 3.095 ;
        RECT  0.150 0.820 0.185 3.095 ;
    END
END MX3X4

MACRO MX3X2
    CLASS CORE ;
    FOREIGN MX3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 0.645 7.695 3.215 ;
        RECT  7.435 0.645 7.535 0.905 ;
        RECT  7.405 2.275 7.535 3.215 ;
        END
        ANTENNADIFFAREA     0.7140 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.960 6.785 2.220 ;
        RECT  6.525 1.960 6.775 2.400 ;
        RECT  6.320 2.240 6.525 2.400 ;
        RECT  6.160 2.240 6.320 2.765 ;
        RECT  4.970 2.605 6.160 2.765 ;
        RECT  4.710 2.505 4.970 2.765 ;
        END
        ANTENNAGATEAREA     0.3432 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.210 2.540 3.260 2.800 ;
        RECT  3.095 2.530 3.210 2.800 ;
        RECT  2.885 2.520 3.095 2.810 ;
        RECT  1.705 2.530 2.885 2.690 ;
        RECT  2.375 0.505 2.635 0.765 ;
        RECT  2.120 0.605 2.375 0.765 ;
        RECT  1.960 0.605 2.120 0.795 ;
        RECT  0.875 0.635 1.960 0.795 ;
        RECT  1.445 2.530 1.705 2.750 ;
        RECT  1.145 2.530 1.445 2.690 ;
        RECT  1.145 1.465 1.185 1.625 ;
        RECT  0.985 1.465 1.145 2.690 ;
        RECT  0.875 1.465 0.985 1.625 ;
        RECT  0.715 0.635 0.875 1.625 ;
        RECT  0.585 1.105 0.715 1.625 ;
        END
        ANTENNAGATEAREA     0.3835 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 1.895 0.795 2.460 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.760 1.290 2.185 1.625 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.290 4.475 1.810 ;
        RECT  4.080 1.550 4.265 1.810 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 -0.250 7.820 0.250 ;
        RECT  6.925 -0.250 7.185 0.885 ;
        RECT  4.485 -0.250 6.925 0.250 ;
        RECT  4.225 -0.250 4.485 0.405 ;
        RECT  1.770 -0.250 4.225 0.250 ;
        RECT  1.510 -0.250 1.770 0.405 ;
        RECT  0.935 -0.250 1.510 0.250 ;
        RECT  0.675 -0.250 0.935 0.450 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.155 3.440 7.820 3.940 ;
        RECT  6.895 2.955 7.155 3.940 ;
        RECT  4.590 3.440 6.895 3.940 ;
        RECT  4.330 3.285 4.590 3.940 ;
        RECT  1.930 3.440 4.330 3.940 ;
        RECT  1.670 3.285 1.930 3.940 ;
        RECT  0.985 3.440 1.670 3.940 ;
        RECT  0.725 3.270 0.985 3.940 ;
        RECT  0.000 3.440 0.725 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.195 1.115 7.355 2.085 ;
        RECT  6.675 1.115 7.195 1.275 ;
        RECT  7.155 1.925 7.195 2.085 ;
        RECT  6.995 1.925 7.155 2.765 ;
        RECT  6.755 1.475 7.015 1.735 ;
        RECT  6.675 2.605 6.995 2.765 ;
        RECT  6.165 1.505 6.755 1.675 ;
        RECT  6.415 0.675 6.675 1.275 ;
        RECT  6.515 2.605 6.675 3.105 ;
        RECT  3.880 2.945 6.515 3.105 ;
        RECT  5.960 0.675 6.165 1.675 ;
        RECT  5.905 0.675 5.960 2.425 ;
        RECT  5.800 1.515 5.905 2.425 ;
        RECT  5.555 0.590 5.655 1.230 ;
        RECT  5.395 0.590 5.555 2.320 ;
        RECT  3.415 0.590 5.395 0.750 ;
        RECT  5.240 2.060 5.395 2.320 ;
        RECT  5.065 1.275 5.205 1.535 ;
        RECT  4.990 0.955 5.065 1.535 ;
        RECT  4.830 0.955 4.990 2.215 ;
        RECT  4.805 0.955 4.830 1.115 ;
        RECT  4.730 1.955 4.830 2.215 ;
        RECT  3.850 2.075 4.040 2.675 ;
        RECT  3.850 0.975 3.925 1.235 ;
        RECT  3.720 2.945 3.880 3.220 ;
        RECT  3.780 0.975 3.850 2.675 ;
        RECT  3.690 0.975 3.780 2.455 ;
        RECT  2.360 3.060 3.720 3.220 ;
        RECT  3.665 0.975 3.690 1.235 ;
        RECT  3.360 2.050 3.460 2.310 ;
        RECT  3.360 0.590 3.415 1.190 ;
        RECT  3.200 0.590 3.360 2.310 ;
        RECT  3.155 0.590 3.200 1.190 ;
        RECT  2.810 0.945 2.970 2.340 ;
        RECT  2.300 0.945 2.810 1.105 ;
        RECT  2.220 2.180 2.810 2.340 ;
        RECT  2.455 1.540 2.615 2.000 ;
        RECT  1.540 1.840 2.455 2.000 ;
        RECT  2.200 2.930 2.360 3.220 ;
        RECT  0.335 2.930 2.200 3.090 ;
        RECT  1.380 1.080 1.540 2.250 ;
        RECT  1.355 1.080 1.380 1.240 ;
        RECT  1.325 1.990 1.380 2.250 ;
        RECT  1.095 0.980 1.355 1.240 ;
        RECT  0.335 0.525 0.385 1.125 ;
        RECT  0.175 0.525 0.335 3.215 ;
        RECT  0.125 0.525 0.175 1.125 ;
    END
END MX3X2

MACRO MX3X1
    CLASS CORE ;
    FOREIGN MX3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.615 0.595 6.775 2.645 ;
        RECT  6.515 0.595 6.615 0.855 ;
        RECT  6.515 1.925 6.615 2.645 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 0.470 4.700 0.720 ;
        RECT  4.265 0.470 4.475 0.760 ;
        RECT  4.180 0.470 4.265 0.720 ;
        END
        ANTENNAGATEAREA     0.1885 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.675 2.930 1.255 3.220 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.635 0.395 1.895 ;
        RECT  0.135 1.635 0.335 2.400 ;
        RECT  0.125 1.895 0.135 2.400 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.315 1.945 1.575 ;
        RECT  1.505 1.290 1.715 1.580 ;
        RECT  1.430 1.315 1.505 1.575 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.640 1.620 4.015 1.990 ;
        RECT  3.480 1.475 3.640 1.990 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.225 -0.250 6.900 0.250 ;
        RECT  5.965 -0.250 6.225 0.405 ;
        RECT  3.855 -0.250 5.965 0.250 ;
        RECT  3.595 -0.250 3.855 1.020 ;
        RECT  1.755 -0.250 3.595 0.250 ;
        RECT  3.555 0.760 3.595 1.020 ;
        RECT  1.495 -0.250 1.755 1.045 ;
        RECT  0.385 -0.250 1.495 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.375 3.440 6.900 3.940 ;
        RECT  6.115 3.285 6.375 3.940 ;
        RECT  3.900 3.440 6.115 3.940 ;
        RECT  3.640 3.285 3.900 3.940 ;
        RECT  1.600 3.440 3.640 3.940 ;
        RECT  1.440 2.915 1.600 3.940 ;
        RECT  0.385 3.440 1.440 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.330 1.070 6.420 1.330 ;
        RECT  6.170 0.690 6.330 1.330 ;
        RECT  5.430 0.690 6.170 0.850 ;
        RECT  6.160 1.070 6.170 1.330 ;
        RECT  5.865 1.125 5.970 1.385 ;
        RECT  5.765 1.125 5.865 2.640 ;
        RECT  5.705 1.125 5.765 3.100 ;
        RECT  5.605 2.380 5.705 3.100 ;
        RECT  2.255 2.940 5.605 3.100 ;
        RECT  5.380 0.690 5.430 1.240 ;
        RECT  5.270 0.690 5.380 2.665 ;
        RECT  5.220 0.980 5.270 2.665 ;
        RECT  5.170 0.980 5.220 1.240 ;
        RECT  5.095 2.405 5.220 2.665 ;
        RECT  4.845 0.945 4.965 2.125 ;
        RECT  4.805 0.945 4.845 2.760 ;
        RECT  4.660 0.945 4.805 1.205 ;
        RECT  4.685 1.965 4.805 2.760 ;
        RECT  2.960 2.600 4.685 2.760 ;
        RECT  4.460 1.510 4.600 1.770 ;
        RECT  4.300 0.960 4.460 2.415 ;
        RECT  4.150 0.960 4.300 1.220 ;
        RECT  4.075 2.255 4.300 2.415 ;
        RECT  3.140 0.755 3.300 2.415 ;
        RECT  3.040 0.755 3.140 0.915 ;
        RECT  2.800 1.100 2.960 2.760 ;
        RECT  2.775 1.100 2.800 1.260 ;
        RECT  2.515 2.600 2.800 2.760 ;
        RECT  2.615 0.755 2.775 1.260 ;
        RECT  2.460 1.440 2.620 2.390 ;
        RECT  2.515 0.755 2.615 1.015 ;
        RECT  2.315 1.440 2.460 1.600 ;
        RECT  1.930 2.230 2.460 2.390 ;
        RECT  2.155 0.780 2.315 1.600 ;
        RECT  2.120 1.780 2.280 2.045 ;
        RECT  2.095 2.570 2.255 3.100 ;
        RECT  2.005 0.780 2.155 1.040 ;
        RECT  1.185 1.885 2.120 2.045 ;
        RECT  0.785 2.570 2.095 2.730 ;
        RECT  1.025 0.520 1.185 2.215 ;
        RECT  0.925 0.520 1.025 0.780 ;
        RECT  0.915 1.955 1.025 2.215 ;
        RECT  0.735 1.030 0.785 1.290 ;
        RECT  0.735 2.470 0.785 2.730 ;
        RECT  0.575 1.030 0.735 2.730 ;
        RECT  0.525 1.030 0.575 1.290 ;
        RECT  0.525 2.470 0.575 2.730 ;
    END
END MX3X1

MACRO MX3XL
    CLASS CORE ;
    FOREIGN MX3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.765 0.430 5.875 2.810 ;
        RECT  5.715 0.430 5.765 2.885 ;
        RECT  5.580 0.430 5.715 0.590 ;
        RECT  5.645 1.925 5.715 2.885 ;
        RECT  5.505 2.625 5.645 2.885 ;
        END
        ANTENNADIFFAREA     0.3370 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 0.435 4.660 0.595 ;
        RECT  3.805 0.435 4.015 0.760 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 2.910 0.520 3.225 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 2.110 5.395 2.400 ;
        RECT  4.900 2.110 5.185 2.370 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.735 1.290 1.255 1.600 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.475 3.120 1.990 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.330 -0.250 5.980 0.250 ;
        RECT  5.070 -0.250 5.330 0.405 ;
        RECT  2.990 -0.250 5.070 0.250 ;
        RECT  2.730 -0.250 2.990 0.405 ;
        RECT  0.955 -0.250 2.730 0.250 ;
        RECT  0.695 -0.250 0.955 1.080 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.350 3.440 5.980 3.940 ;
        RECT  5.090 3.285 5.350 3.940 ;
        RECT  3.140 3.440 5.090 3.940 ;
        RECT  2.880 3.285 3.140 3.940 ;
        RECT  0.960 3.440 2.880 3.940 ;
        RECT  0.700 2.740 0.960 3.940 ;
        RECT  0.000 3.440 0.700 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.375 1.000 5.535 1.515 ;
        RECT  4.495 1.000 5.375 1.160 ;
        RECT  4.720 1.340 4.890 1.600 ;
        RECT  4.720 2.665 4.770 2.925 ;
        RECT  4.560 1.340 4.720 2.925 ;
        RECT  4.510 2.665 4.560 2.925 ;
        RECT  4.380 0.810 4.495 1.160 ;
        RECT  4.220 0.810 4.380 2.410 ;
        RECT  4.205 2.250 4.220 2.410 ;
        RECT  4.045 2.250 4.205 3.040 ;
        RECT  3.880 1.025 4.040 2.070 ;
        RECT  3.690 1.025 3.880 1.285 ;
        RECT  3.865 1.910 3.880 2.070 ;
        RECT  3.725 1.910 3.865 2.760 ;
        RECT  3.705 1.910 3.725 2.925 ;
        RECT  3.465 2.600 3.705 2.925 ;
        RECT  3.480 1.470 3.690 1.730 ;
        RECT  3.480 0.515 3.580 0.775 ;
        RECT  3.480 2.155 3.520 2.415 ;
        RECT  3.320 0.515 3.480 2.415 ;
        RECT  2.130 2.600 3.465 2.760 ;
        RECT  2.335 0.820 2.495 2.415 ;
        RECT  1.970 0.820 2.130 2.760 ;
        RECT  1.775 0.820 1.970 1.080 ;
        RECT  1.930 2.565 1.970 2.760 ;
        RECT  1.670 2.565 1.930 2.825 ;
        RECT  1.630 1.435 1.790 2.385 ;
        RECT  1.595 1.435 1.630 1.595 ;
        RECT  1.390 2.225 1.630 2.385 ;
        RECT  1.435 0.820 1.595 1.595 ;
        RECT  1.290 1.780 1.450 2.040 ;
        RECT  1.265 0.820 1.435 1.080 ;
        RECT  1.130 2.225 1.390 2.485 ;
        RECT  0.385 1.780 1.290 1.940 ;
        RECT  0.225 0.820 0.385 2.415 ;
        RECT  0.125 0.820 0.225 1.080 ;
        RECT  0.125 2.155 0.225 2.415 ;
    END
END MX3XL

MACRO MXI4X4
    CLASS CORE ;
    FOREIGN MXI4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.535 0.630 9.600 2.605 ;
        RECT  9.485 0.630 9.535 2.810 ;
        RECT  9.400 0.630 9.485 2.975 ;
        RECT  9.225 0.630 9.400 0.890 ;
        RECT  9.225 2.035 9.400 2.975 ;
        END
        ANTENNADIFFAREA     0.8592 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.290 7.815 1.935 ;
        END
        ANTENNAGATEAREA     0.3536 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.700 2.715 2.140 ;
        END
        ANTENNAGATEAREA     0.5382 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.245 1.290 3.555 1.740 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.095 1.130 5.395 1.670 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 1.265 2.245 1.665 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.585 0.395 1.845 ;
        RECT  0.130 1.585 0.335 2.810 ;
        RECT  0.125 1.925 0.130 2.810 ;
        END
        ANTENNAGATEAREA     0.1950 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.945 -0.250 10.120 0.250 ;
        RECT  9.785 -0.250 9.945 1.095 ;
        RECT  8.835 -0.250 9.785 0.250 ;
        RECT  8.575 -0.250 8.835 0.405 ;
        RECT  7.885 -0.250 8.575 0.250 ;
        RECT  7.625 -0.250 7.885 0.405 ;
        RECT  5.415 -0.250 7.625 0.250 ;
        RECT  5.155 -0.250 5.415 0.950 ;
        RECT  3.300 -0.250 5.155 0.250 ;
        RECT  3.040 -0.250 3.300 0.575 ;
        RECT  2.425 -0.250 3.040 0.250 ;
        RECT  2.165 -0.250 2.425 1.085 ;
        RECT  0.385 -0.250 2.165 0.250 ;
        RECT  0.125 -0.250 0.385 0.865 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.995 3.440 10.120 3.940 ;
        RECT  9.945 2.935 9.995 3.940 ;
        RECT  9.785 2.250 9.945 3.940 ;
        RECT  9.735 2.935 9.785 3.940 ;
        RECT  8.945 3.440 9.735 3.940 ;
        RECT  8.685 3.285 8.945 3.940 ;
        RECT  7.980 3.440 8.685 3.940 ;
        RECT  7.720 3.285 7.980 3.940 ;
        RECT  5.415 3.440 7.720 3.940 ;
        RECT  5.155 3.285 5.415 3.940 ;
        RECT  3.265 3.440 5.155 3.940 ;
        RECT  3.005 3.110 3.265 3.940 ;
        RECT  2.485 3.440 3.005 3.940 ;
        RECT  2.225 3.110 2.485 3.940 ;
        RECT  0.385 3.440 2.225 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.060 1.070 9.220 1.775 ;
        RECT  8.775 1.070 9.060 1.230 ;
        RECT  8.700 1.510 8.860 3.105 ;
        RECT  8.615 0.585 8.775 1.230 ;
        RECT  8.695 1.510 8.700 1.670 ;
        RECT  3.605 2.945 8.700 3.105 ;
        RECT  8.435 1.410 8.695 1.670 ;
        RECT  6.460 0.585 8.615 0.745 ;
        RECT  8.360 1.850 8.520 2.765 ;
        RECT  8.175 0.965 8.435 1.225 ;
        RECT  8.155 1.850 8.360 2.010 ;
        RECT  6.800 2.605 8.360 2.765 ;
        RECT  8.155 1.065 8.175 1.225 ;
        RECT  7.995 1.065 8.155 2.010 ;
        RECT  7.270 2.160 7.595 2.420 ;
        RECT  7.270 0.925 7.485 1.085 ;
        RECT  7.110 0.925 7.270 2.420 ;
        RECT  6.980 1.405 7.110 1.565 ;
        RECT  6.800 0.925 6.925 1.185 ;
        RECT  6.640 0.925 6.800 2.765 ;
        RECT  6.300 0.585 6.460 2.765 ;
        RECT  6.255 0.585 6.300 1.065 ;
        RECT  6.255 2.165 6.300 2.765 ;
        RECT  5.915 0.645 6.075 2.735 ;
        RECT  5.695 0.645 5.915 1.245 ;
        RECT  5.695 2.235 5.915 2.735 ;
        RECT  5.575 1.670 5.735 2.055 ;
        RECT  5.255 1.895 5.575 2.055 ;
        RECT  5.095 1.895 5.255 2.765 ;
        RECT  4.575 2.605 5.095 2.765 ;
        RECT  4.755 0.745 4.915 2.425 ;
        RECT  4.610 0.745 4.755 0.905 ;
        RECT  4.415 1.085 4.575 2.765 ;
        RECT  4.360 1.085 4.415 1.245 ;
        RECT  4.055 2.605 4.415 2.765 ;
        RECT  4.200 0.850 4.360 1.245 ;
        RECT  4.075 1.435 4.235 2.425 ;
        RECT  4.100 0.850 4.200 1.110 ;
        RECT  3.895 1.435 4.075 1.595 ;
        RECT  3.805 2.265 4.075 2.425 ;
        RECT  3.735 0.850 3.895 1.595 ;
        RECT  3.735 1.775 3.895 2.085 ;
        RECT  3.545 2.265 3.805 2.525 ;
        RECT  3.590 0.850 3.735 1.110 ;
        RECT  3.065 1.925 3.735 2.085 ;
        RECT  3.445 2.770 3.605 3.105 ;
        RECT  1.345 2.770 3.445 2.930 ;
        RECT  2.935 1.015 3.065 2.480 ;
        RECT  2.905 0.945 2.935 2.480 ;
        RECT  2.675 0.945 2.905 1.205 ;
        RECT  2.895 2.320 2.905 2.480 ;
        RECT  2.635 2.320 2.895 2.580 ;
        RECT  2.200 2.320 2.635 2.480 ;
        RECT  2.040 1.845 2.200 2.480 ;
        RECT  1.755 1.845 2.040 2.005 ;
        RECT  1.745 0.815 1.915 1.075 ;
        RECT  1.805 2.325 1.855 2.585 ;
        RECT  1.595 2.185 1.805 2.585 ;
        RECT  1.595 1.675 1.755 2.005 ;
        RECT  1.585 0.815 1.745 1.495 ;
        RECT  1.415 2.185 1.595 2.345 ;
        RECT  1.415 1.335 1.585 1.495 ;
        RECT  1.255 1.335 1.415 2.345 ;
        RECT  1.145 0.895 1.405 1.155 ;
        RECT  1.075 2.525 1.345 2.930 ;
        RECT  1.075 0.995 1.145 1.155 ;
        RECT  0.915 0.995 1.075 2.930 ;
        RECT  0.735 0.655 0.895 0.815 ;
        RECT  0.575 0.655 0.735 2.655 ;
    END
END MXI4X4

MACRO MXI4X2
    CLASS CORE ;
    FOREIGN MXI4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.355 0.695 9.535 3.045 ;
        RECT  9.275 0.495 9.355 3.045 ;
        RECT  9.095 0.495 9.275 1.095 ;
        END
        ANTENNADIFFAREA     0.7272 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.445 1.290 7.695 1.890 ;
        END
        ANTENNAGATEAREA     0.2951 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.420 1.315 2.635 2.000 ;
        RECT  2.385 1.740 2.420 2.000 ;
        END
        ANTENNAGATEAREA     0.4524 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.290 3.555 1.580 ;
        RECT  3.345 1.290 3.500 1.745 ;
        RECT  3.195 1.295 3.345 1.745 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.095 1.280 5.475 1.615 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 1.185 2.205 1.660 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.135 1.585 0.395 2.150 ;
        RECT  0.125 1.700 0.135 2.150 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.815 -0.250 9.660 0.250 ;
        RECT  8.555 -0.250 8.815 1.090 ;
        RECT  7.435 -0.250 8.555 0.250 ;
        RECT  7.175 -0.250 7.435 0.405 ;
        RECT  5.385 -0.250 7.175 0.250 ;
        RECT  5.125 -0.250 5.385 0.875 ;
        RECT  3.395 -0.250 5.125 0.250 ;
        RECT  3.135 -0.250 3.395 0.575 ;
        RECT  2.375 -0.250 3.135 0.250 ;
        RECT  2.115 -0.250 2.375 1.005 ;
        RECT  0.385 -0.250 2.115 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.965 3.440 9.660 3.940 ;
        RECT  8.965 2.215 8.970 3.155 ;
        RECT  8.785 2.215 8.965 3.940 ;
        RECT  8.705 3.285 8.785 3.940 ;
        RECT  7.765 3.440 8.705 3.940 ;
        RECT  7.505 3.285 7.765 3.940 ;
        RECT  5.365 3.440 7.505 3.940 ;
        RECT  5.105 3.285 5.365 3.940 ;
        RECT  3.265 3.440 5.105 3.940 ;
        RECT  3.005 3.110 3.265 3.940 ;
        RECT  2.485 3.440 3.005 3.940 ;
        RECT  2.225 3.110 2.485 3.940 ;
        RECT  0.385 3.440 2.225 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.935 1.280 9.095 1.665 ;
        RECT  8.375 1.280 8.935 1.440 ;
        RECT  8.445 1.625 8.605 3.105 ;
        RECT  8.260 1.625 8.445 1.785 ;
        RECT  7.320 2.945 8.445 3.105 ;
        RECT  8.215 0.585 8.375 1.440 ;
        RECT  8.035 2.165 8.265 2.765 ;
        RECT  6.415 0.585 8.215 0.745 ;
        RECT  7.875 1.035 8.035 2.765 ;
        RECT  6.975 2.605 7.875 2.765 ;
        RECT  7.265 0.950 7.485 1.110 ;
        RECT  7.265 2.210 7.375 2.370 ;
        RECT  7.160 2.945 7.320 3.220 ;
        RECT  7.105 0.950 7.265 2.370 ;
        RECT  5.925 3.060 7.160 3.220 ;
        RECT  6.935 1.405 7.105 1.665 ;
        RECT  6.755 2.605 6.975 2.880 ;
        RECT  6.765 0.925 6.925 1.185 ;
        RECT  6.755 0.980 6.765 1.185 ;
        RECT  6.595 0.980 6.755 2.880 ;
        RECT  6.365 0.585 6.415 1.065 ;
        RECT  6.365 2.165 6.415 2.765 ;
        RECT  6.205 0.585 6.365 2.765 ;
        RECT  5.795 0.565 5.955 2.735 ;
        RECT  5.765 2.945 5.925 3.220 ;
        RECT  5.695 0.565 5.795 1.165 ;
        RECT  5.695 2.235 5.795 2.735 ;
        RECT  3.605 2.945 5.765 3.105 ;
        RECT  5.515 1.795 5.615 2.055 ;
        RECT  5.355 1.795 5.515 2.765 ;
        RECT  4.575 2.605 5.355 2.765 ;
        RECT  4.755 0.665 4.915 2.425 ;
        RECT  4.615 0.665 4.755 0.825 ;
        RECT  4.415 1.005 4.575 2.765 ;
        RECT  4.335 1.005 4.415 1.165 ;
        RECT  4.055 2.605 4.415 2.765 ;
        RECT  4.075 0.905 4.335 1.165 ;
        RECT  4.075 1.355 4.235 2.425 ;
        RECT  3.895 1.355 4.075 1.515 ;
        RECT  3.805 2.265 4.075 2.425 ;
        RECT  3.735 0.950 3.895 1.515 ;
        RECT  3.735 1.695 3.895 2.085 ;
        RECT  3.545 2.265 3.805 2.525 ;
        RECT  3.565 0.950 3.735 1.110 ;
        RECT  2.975 1.925 3.735 2.085 ;
        RECT  3.445 2.770 3.605 3.105 ;
        RECT  1.295 2.770 3.445 2.930 ;
        RECT  2.815 0.825 2.975 2.340 ;
        RECT  2.625 0.825 2.815 1.085 ;
        RECT  2.145 2.180 2.815 2.340 ;
        RECT  1.985 1.840 2.145 2.340 ;
        RECT  1.755 1.840 1.985 2.000 ;
        RECT  1.735 0.745 1.835 1.005 ;
        RECT  1.545 2.180 1.805 2.585 ;
        RECT  1.595 1.740 1.755 2.000 ;
        RECT  1.575 0.745 1.735 1.505 ;
        RECT  1.415 1.345 1.575 1.505 ;
        RECT  1.415 2.180 1.545 2.340 ;
        RECT  1.255 1.345 1.415 2.340 ;
        RECT  1.075 0.885 1.325 1.145 ;
        RECT  1.075 2.570 1.295 2.930 ;
        RECT  1.065 0.885 1.075 2.930 ;
        RECT  0.915 0.980 1.065 2.930 ;
        RECT  0.575 1.035 0.735 2.405 ;
    END
END MXI4X2

MACRO MXI4X1
    CLASS CORE ;
    FOREIGN MXI4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.455 0.545 8.615 2.400 ;
        RECT  8.355 0.545 8.455 0.805 ;
        RECT  8.405 1.925 8.455 2.400 ;
        RECT  7.995 2.175 8.405 2.400 ;
        RECT  7.735 2.175 7.995 2.435 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.595 7.815 1.990 ;
        RECT  7.480 1.595 7.485 1.855 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 1.700 2.635 2.220 ;
        RECT  2.340 2.060 2.355 2.220 ;
        END
        ANTENNAGATEAREA     0.2275 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.290 4.015 1.580 ;
        RECT  3.755 1.340 3.805 1.580 ;
        RECT  3.495 1.340 3.755 1.600 ;
        END
        ANTENNAGATEAREA     0.0793 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 1.290 5.395 1.580 ;
        RECT  5.035 1.355 5.185 1.580 ;
        RECT  4.875 1.355 5.035 1.720 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.185 2.280 1.520 ;
        RECT  1.945 1.185 2.175 1.580 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.845 0.335 2.810 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.075 -0.250 8.740 0.250 ;
        RECT  7.815 -0.250 8.075 0.405 ;
        RECT  7.220 -0.250 7.815 0.250 ;
        RECT  6.960 -0.250 7.220 0.625 ;
        RECT  5.185 -0.250 6.960 0.250 ;
        RECT  4.925 -0.250 5.185 0.795 ;
        RECT  2.920 -0.250 4.925 0.250 ;
        RECT  2.760 -0.250 2.920 0.875 ;
        RECT  2.390 -0.250 2.760 0.250 ;
        RECT  2.130 -0.250 2.390 1.005 ;
        RECT  0.385 -0.250 2.130 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.535 3.440 8.740 3.940 ;
        RECT  8.275 2.605 8.535 3.940 ;
        RECT  7.265 3.440 8.275 3.940 ;
        RECT  7.105 2.955 7.265 3.940 ;
        RECT  5.210 3.440 7.105 3.940 ;
        RECT  4.950 3.285 5.210 3.940 ;
        RECT  3.140 3.440 4.950 3.940 ;
        RECT  2.880 3.115 3.140 3.940 ;
        RECT  2.205 3.440 2.880 3.940 ;
        RECT  1.945 3.115 2.205 3.940 ;
        RECT  0.385 3.440 1.945 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.175 0.985 8.275 1.245 ;
        RECT  8.015 0.805 8.175 1.245 ;
        RECT  6.125 0.805 8.015 0.965 ;
        RECT  7.785 2.970 7.885 3.230 ;
        RECT  7.295 1.175 7.795 1.335 ;
        RECT  7.625 2.615 7.785 3.230 ;
        RECT  7.295 2.615 7.625 2.775 ;
        RECT  7.135 1.175 7.295 2.775 ;
        RECT  6.595 1.655 7.135 1.915 ;
        RECT  6.765 2.135 6.925 3.105 ;
        RECT  4.515 2.945 6.765 3.105 ;
        RECT  6.415 1.180 6.715 1.340 ;
        RECT  6.425 2.155 6.585 2.765 ;
        RECT  6.415 2.155 6.425 2.315 ;
        RECT  6.255 1.180 6.415 2.315 ;
        RECT  6.075 0.805 6.125 0.970 ;
        RECT  5.915 0.805 6.075 2.755 ;
        RECT  5.575 1.370 5.735 2.640 ;
        RECT  5.350 2.380 5.575 2.640 ;
        RECT  5.050 1.940 5.310 2.200 ;
        RECT  5.035 2.040 5.050 2.200 ;
        RECT  4.875 2.040 5.035 2.760 ;
        RECT  4.190 2.600 4.875 2.760 ;
        RECT  4.535 1.090 4.695 2.365 ;
        RECT  4.370 2.105 4.535 2.365 ;
        RECT  4.355 2.945 4.515 3.150 ;
        RECT  4.195 0.950 4.355 1.920 ;
        RECT  3.705 2.990 4.355 3.150 ;
        RECT  4.110 0.950 4.195 1.110 ;
        RECT  4.190 1.760 4.195 1.920 ;
        RECT  4.095 1.760 4.190 2.760 ;
        RECT  3.850 0.850 4.110 1.110 ;
        RECT  4.030 1.760 4.095 2.810 ;
        RECT  3.935 2.550 4.030 2.810 ;
        RECT  3.755 1.820 3.780 2.080 ;
        RECT  3.595 1.820 3.755 2.595 ;
        RECT  3.545 2.775 3.705 3.150 ;
        RECT  2.975 2.435 3.595 2.595 ;
        RECT  1.325 2.775 3.545 2.935 ;
        RECT  3.315 0.685 3.540 0.945 ;
        RECT  3.315 2.095 3.415 2.255 ;
        RECT  3.155 0.685 3.315 2.255 ;
        RECT  2.815 1.125 2.975 2.595 ;
        RECT  2.710 1.125 2.815 1.385 ;
        RECT  2.075 2.435 2.815 2.595 ;
        RECT  1.915 1.795 2.075 2.595 ;
        RECT  1.760 1.795 1.915 1.955 ;
        RECT  1.600 1.695 1.760 1.955 ;
        RECT  1.590 1.005 1.750 1.290 ;
        RECT  1.475 2.260 1.735 2.520 ;
        RECT  1.420 1.130 1.590 1.290 ;
        RECT  1.420 2.260 1.475 2.420 ;
        RECT  1.260 1.130 1.420 2.420 ;
        RECT  1.080 2.775 1.325 3.140 ;
        RECT  1.080 0.505 1.220 0.765 ;
        RECT  1.065 0.505 1.080 3.140 ;
        RECT  0.960 0.505 1.065 2.935 ;
        RECT  0.920 0.525 0.960 2.935 ;
        RECT  0.675 1.035 0.740 1.295 ;
        RECT  0.675 2.260 0.735 2.520 ;
        RECT  0.515 1.035 0.675 2.520 ;
    END
END MXI4X1

MACRO MXI4XL
    CLASS CORE ;
    FOREIGN MXI4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.455 0.615 8.615 2.400 ;
        RECT  8.430 0.615 8.455 0.945 ;
        RECT  8.405 1.925 8.455 2.400 ;
        RECT  8.355 0.615 8.430 0.875 ;
        RECT  7.705 2.170 8.405 2.400 ;
        END
        ANTENNADIFFAREA     0.2597 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.830 1.700 8.155 1.990 ;
        RECT  7.570 1.595 7.830 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.390 1.565 2.635 2.220 ;
        RECT  2.340 2.060 2.390 2.220 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.290 4.015 1.580 ;
        RECT  3.755 1.335 3.805 1.580 ;
        RECT  3.495 1.335 3.755 1.595 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 1.290 5.395 1.580 ;
        RECT  5.035 1.355 5.185 1.580 ;
        RECT  4.875 1.355 5.035 1.720 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 1.290 2.210 1.815 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.845 0.335 2.810 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.035 -0.250 8.740 0.250 ;
        RECT  7.775 -0.250 8.035 0.405 ;
        RECT  7.220 -0.250 7.775 0.250 ;
        RECT  6.960 -0.250 7.220 0.625 ;
        RECT  5.185 -0.250 6.960 0.250 ;
        RECT  4.925 -0.250 5.185 0.795 ;
        RECT  2.920 -0.250 4.925 0.250 ;
        RECT  2.760 -0.250 2.920 0.875 ;
        RECT  2.395 -0.250 2.760 0.250 ;
        RECT  2.135 -0.250 2.395 1.110 ;
        RECT  0.385 -0.250 2.135 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.535 3.440 8.740 3.940 ;
        RECT  8.275 2.605 8.535 3.940 ;
        RECT  7.405 3.440 8.275 3.940 ;
        RECT  7.245 2.955 7.405 3.940 ;
        RECT  5.160 3.440 7.245 3.940 ;
        RECT  4.900 3.285 5.160 3.940 ;
        RECT  3.135 3.440 4.900 3.940 ;
        RECT  2.875 3.115 3.135 3.940 ;
        RECT  2.185 3.440 2.875 3.940 ;
        RECT  1.925 3.115 2.185 3.940 ;
        RECT  0.385 3.440 1.925 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.145 1.060 8.245 1.320 ;
        RECT  7.985 0.805 8.145 1.320 ;
        RECT  7.925 2.970 8.025 3.230 ;
        RECT  6.205 0.805 7.985 0.965 ;
        RECT  7.765 2.615 7.925 3.230 ;
        RECT  7.390 1.175 7.795 1.335 ;
        RECT  7.390 2.615 7.765 2.775 ;
        RECT  7.230 1.175 7.390 2.775 ;
        RECT  6.595 1.655 7.230 1.925 ;
        RECT  7.020 2.135 7.050 2.410 ;
        RECT  6.860 2.135 7.020 3.105 ;
        RECT  4.535 2.945 6.860 3.105 ;
        RECT  6.675 1.175 6.725 1.335 ;
        RECT  6.520 2.105 6.680 2.615 ;
        RECT  6.465 1.175 6.675 1.340 ;
        RECT  6.415 2.105 6.520 2.265 ;
        RECT  6.415 1.180 6.465 1.340 ;
        RECT  6.255 1.180 6.415 2.265 ;
        RECT  6.075 0.695 6.205 0.965 ;
        RECT  6.075 2.450 6.110 2.715 ;
        RECT  5.915 0.695 6.075 2.715 ;
        RECT  5.575 1.205 5.735 2.640 ;
        RECT  5.330 2.380 5.575 2.640 ;
        RECT  5.050 1.940 5.310 2.200 ;
        RECT  5.035 2.040 5.050 2.200 ;
        RECT  4.875 2.040 5.035 2.700 ;
        RECT  4.120 2.540 4.875 2.700 ;
        RECT  4.535 1.090 4.695 2.360 ;
        RECT  4.305 2.100 4.535 2.360 ;
        RECT  4.375 2.945 4.535 3.210 ;
        RECT  3.755 3.050 4.375 3.210 ;
        RECT  4.195 0.950 4.355 1.920 ;
        RECT  4.110 0.950 4.195 1.110 ;
        RECT  4.120 1.760 4.195 1.920 ;
        RECT  3.960 1.760 4.120 2.870 ;
        RECT  3.850 0.850 4.110 1.110 ;
        RECT  3.935 2.540 3.960 2.870 ;
        RECT  3.755 1.820 3.780 2.085 ;
        RECT  3.595 1.820 3.755 2.595 ;
        RECT  3.595 2.775 3.755 3.210 ;
        RECT  2.975 2.435 3.595 2.595 ;
        RECT  1.325 2.775 3.595 2.935 ;
        RECT  3.315 0.795 3.540 1.055 ;
        RECT  3.315 2.095 3.415 2.255 ;
        RECT  3.155 0.795 3.315 2.255 ;
        RECT  2.815 1.125 2.975 2.595 ;
        RECT  2.710 1.125 2.815 1.385 ;
        RECT  2.095 2.435 2.815 2.595 ;
        RECT  1.935 1.995 2.095 2.595 ;
        RECT  1.715 1.995 1.935 2.155 ;
        RECT  1.615 1.035 1.775 1.665 ;
        RECT  1.495 2.335 1.755 2.595 ;
        RECT  1.555 1.845 1.715 2.155 ;
        RECT  1.375 1.505 1.615 1.665 ;
        RECT  1.375 2.335 1.495 2.495 ;
        RECT  1.215 1.505 1.375 2.495 ;
        RECT  1.065 2.775 1.325 3.140 ;
        RECT  1.035 1.035 1.255 1.295 ;
        RECT  1.035 2.775 1.065 2.935 ;
        RECT  0.875 1.035 1.035 2.935 ;
        RECT  0.845 0.525 0.895 0.785 ;
        RECT  0.695 0.525 0.845 0.815 ;
        RECT  0.635 0.525 0.695 2.985 ;
        RECT  0.535 0.655 0.635 2.985 ;
    END
END MXI4XL

MACRO MXI2X8
    CLASS CORE ;
    FOREIGN MXI2X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.020 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.830 0.695 16.895 2.810 ;
        RECT  16.760 0.585 16.830 2.810 ;
        RECT  16.540 0.585 16.760 3.105 ;
        RECT  13.635 0.585 16.540 0.875 ;
        RECT  16.225 2.110 16.540 3.105 ;
        RECT  11.740 2.705 16.225 3.105 ;
        RECT  3.095 0.585 13.635 0.845 ;
        RECT  2.890 2.775 11.740 3.105 ;
        END
        ANTENNADIFFAREA     5.8484 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.520 1.415 15.780 1.595 ;
        RECT  14.850 1.415 15.520 1.575 ;
        RECT  14.690 1.415 14.850 1.930 ;
        RECT  14.080 1.770 14.690 1.930 ;
        RECT  13.920 1.415 14.080 1.930 ;
        RECT  13.160 1.415 13.920 1.575 ;
        RECT  13.000 1.415 13.160 1.930 ;
        RECT  12.380 1.770 13.000 1.930 ;
        RECT  12.220 1.365 12.380 1.930 ;
        RECT  12.120 1.365 12.220 1.625 ;
        RECT  11.510 1.365 12.120 1.525 ;
        RECT  11.350 1.365 11.510 1.930 ;
        RECT  10.830 1.770 11.350 1.930 ;
        RECT  10.670 1.365 10.830 1.930 ;
        RECT  10.060 1.365 10.670 1.525 ;
        RECT  9.995 1.365 10.060 1.645 ;
        RECT  9.945 1.365 9.995 1.765 ;
        RECT  9.800 1.365 9.945 2.215 ;
        RECT  9.785 1.435 9.800 2.215 ;
        RECT  8.090 2.055 9.785 2.215 ;
        RECT  7.930 1.705 8.090 2.215 ;
        RECT  6.390 2.055 7.930 2.215 ;
        RECT  6.230 1.705 6.390 2.215 ;
        RECT  4.695 2.055 6.230 2.215 ;
        RECT  4.535 1.705 4.695 2.215 ;
        RECT  2.995 2.055 4.535 2.215 ;
        RECT  2.835 1.705 2.995 2.215 ;
        RECT  1.405 2.055 2.835 2.215 ;
        RECT  1.245 1.645 1.405 2.215 ;
        RECT  1.045 1.645 1.245 1.990 ;
        RECT  1.025 1.645 1.045 1.925 ;
        RECT  0.805 1.645 1.025 1.905 ;
        END
        ANTENNAGATEAREA     2.7690 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.160 1.325 16.260 1.585 ;
        RECT  16.000 1.075 16.160 1.585 ;
        RECT  14.510 1.075 16.000 1.235 ;
        RECT  14.350 1.075 14.510 1.590 ;
        RECT  12.820 1.075 14.350 1.235 ;
        RECT  12.660 1.025 12.820 1.590 ;
        RECT  11.170 1.025 12.660 1.185 ;
        RECT  11.010 1.025 11.170 1.590 ;
        RECT  9.580 1.025 11.010 1.185 ;
        RECT  9.420 1.025 9.580 1.605 ;
        RECT  9.325 1.290 9.420 1.605 ;
        RECT  9.320 1.345 9.325 1.605 ;
        END
        ANTENNAGATEAREA     1.9968 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.980 1.515 9.100 1.855 ;
        RECT  8.820 1.025 8.980 1.855 ;
        RECT  7.410 1.025 8.820 1.185 ;
        RECT  7.150 1.025 7.410 1.535 ;
        RECT  5.710 1.025 7.150 1.185 ;
        RECT  5.450 1.025 5.710 1.535 ;
        RECT  4.010 1.025 5.450 1.185 ;
        RECT  3.750 1.025 4.010 1.535 ;
        RECT  2.635 1.025 3.750 1.185 ;
        RECT  2.425 0.880 2.635 1.185 ;
        RECT  2.295 1.025 2.425 1.185 ;
        RECT  2.035 1.025 2.295 1.535 ;
        END
        ANTENNAGATEAREA     1.9968 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.460 -0.250 17.020 0.250 ;
        RECT  16.200 -0.250 16.460 0.405 ;
        RECT  14.760 -0.250 16.200 0.250 ;
        RECT  14.500 -0.250 14.760 0.405 ;
        RECT  13.060 -0.250 14.500 0.250 ;
        RECT  12.800 -0.250 13.060 0.405 ;
        RECT  11.265 -0.250 12.800 0.250 ;
        RECT  11.005 -0.250 11.265 0.405 ;
        RECT  9.350 -0.250 11.005 0.250 ;
        RECT  9.090 -0.250 9.350 0.405 ;
        RECT  7.610 -0.250 9.090 0.250 ;
        RECT  7.350 -0.250 7.610 0.405 ;
        RECT  5.910 -0.250 7.350 0.250 ;
        RECT  5.650 -0.250 5.910 0.405 ;
        RECT  4.205 -0.250 5.650 0.250 ;
        RECT  3.945 -0.250 4.205 0.405 ;
        RECT  2.355 -0.250 3.945 0.250 ;
        RECT  2.220 -0.250 2.355 0.475 ;
        RECT  2.060 -0.250 2.220 0.845 ;
        RECT  1.135 -0.250 2.060 0.250 ;
        RECT  1.960 0.540 2.060 0.845 ;
        RECT  0.875 -0.250 1.135 1.070 ;
        RECT  0.000 -0.250 0.875 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.325 3.440 17.020 3.940 ;
        RECT  16.065 3.285 16.325 3.940 ;
        RECT  14.620 3.440 16.065 3.940 ;
        RECT  14.360 3.285 14.620 3.940 ;
        RECT  12.920 3.440 14.360 3.940 ;
        RECT  12.660 3.285 12.920 3.940 ;
        RECT  11.220 3.440 12.660 3.940 ;
        RECT  10.960 3.285 11.220 3.940 ;
        RECT  9.350 3.440 10.960 3.940 ;
        RECT  9.090 3.285 9.350 3.940 ;
        RECT  7.440 3.440 9.090 3.940 ;
        RECT  7.180 3.285 7.440 3.940 ;
        RECT  5.740 3.440 7.180 3.940 ;
        RECT  5.480 3.285 5.740 3.940 ;
        RECT  4.040 3.440 5.480 3.940 ;
        RECT  3.780 3.285 4.040 3.940 ;
        RECT  2.295 3.440 3.780 3.940 ;
        RECT  2.035 2.935 2.295 3.940 ;
        RECT  1.170 3.440 2.035 3.940 ;
        RECT  0.910 2.895 1.170 3.940 ;
        RECT  0.000 3.440 0.910 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.200 1.755 15.300 1.915 ;
        RECT  15.040 1.755 15.200 2.270 ;
        RECT  13.600 2.110 15.040 2.270 ;
        RECT  13.340 1.755 13.600 2.270 ;
        RECT  11.850 2.110 13.340 2.270 ;
        RECT  11.690 1.705 11.850 2.270 ;
        RECT  10.490 2.110 11.690 2.270 ;
        RECT  10.330 1.705 10.490 2.555 ;
        RECT  1.710 2.395 10.330 2.555 ;
        RECT  8.360 1.365 8.620 1.625 ;
        RECT  7.750 1.365 8.360 1.525 ;
        RECT  7.590 1.365 7.750 1.875 ;
        RECT  6.920 1.715 7.590 1.875 ;
        RECT  6.760 1.365 6.920 1.875 ;
        RECT  6.660 1.365 6.760 1.645 ;
        RECT  6.050 1.365 6.660 1.525 ;
        RECT  5.890 1.365 6.050 1.875 ;
        RECT  5.225 1.715 5.890 1.875 ;
        RECT  5.065 1.365 5.225 1.875 ;
        RECT  4.965 1.365 5.065 1.645 ;
        RECT  4.350 1.365 4.965 1.525 ;
        RECT  4.190 1.365 4.350 1.875 ;
        RECT  3.525 1.715 4.190 1.875 ;
        RECT  3.365 1.365 3.525 1.875 ;
        RECT  3.265 1.365 3.365 1.645 ;
        RECT  2.650 1.365 3.265 1.525 ;
        RECT  2.490 1.365 2.650 1.875 ;
        RECT  1.745 1.715 2.490 1.875 ;
        RECT  1.645 1.305 1.745 1.875 ;
        RECT  1.450 2.395 1.710 3.045 ;
        RECT  1.585 0.615 1.645 1.875 ;
        RECT  1.385 0.615 1.585 1.465 ;
        RECT  0.625 2.395 1.450 2.555 ;
        RECT  0.625 1.305 1.385 1.465 ;
        RECT  0.365 0.695 0.625 3.085 ;
    END
END MXI2X8

MACRO MXI2X6
    CLASS CORE ;
    FOREIGN MXI2X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.220 0.585 12.480 2.810 ;
        RECT  12.110 0.585 12.220 0.945 ;
        RECT  11.925 2.110 12.220 2.810 ;
        RECT  1.115 0.585 12.110 0.845 ;
        RECT  11.585 2.110 11.925 3.105 ;
        RECT  0.945 2.805 11.585 3.105 ;
        END
        ANTENNADIFFAREA     4.3834 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.250 1.365 11.510 1.625 ;
        RECT  10.590 1.365 11.250 1.525 ;
        RECT  10.430 1.365 10.590 2.015 ;
        RECT  9.820 1.855 10.430 2.015 ;
        RECT  9.660 1.365 9.820 2.015 ;
        RECT  9.560 1.365 9.660 1.625 ;
        RECT  8.900 1.365 9.560 1.525 ;
        RECT  8.740 1.365 8.900 1.930 ;
        RECT  8.220 1.770 8.740 1.930 ;
        RECT  8.060 1.365 8.220 1.930 ;
        RECT  7.400 1.365 8.060 1.525 ;
        RECT  7.300 1.365 7.400 1.645 ;
        RECT  7.140 1.365 7.300 2.240 ;
        RECT  6.315 2.080 7.140 2.240 ;
        RECT  5.950 1.635 6.315 2.240 ;
        RECT  4.410 2.080 5.950 2.240 ;
        RECT  4.250 1.705 4.410 2.240 ;
        RECT  2.715 2.080 4.250 2.240 ;
        RECT  2.555 1.705 2.715 2.240 ;
        RECT  1.015 2.080 2.555 2.240 ;
        RECT  0.855 1.705 1.015 2.240 ;
        END
        ANTENNAGATEAREA     2.0124 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.325 12.000 1.585 ;
        RECT  11.740 1.025 11.900 1.585 ;
        RECT  10.250 1.025 11.740 1.185 ;
        RECT  10.005 1.025 10.250 1.675 ;
        RECT  8.560 1.025 10.005 1.185 ;
        RECT  8.400 1.025 8.560 1.590 ;
        RECT  6.920 1.025 8.400 1.185 ;
        RECT  6.760 1.025 6.920 1.605 ;
        RECT  6.660 1.290 6.760 1.605 ;
        RECT  6.565 1.290 6.660 1.580 ;
        END
        ANTENNAGATEAREA     1.4976 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.330 1.395 5.430 1.555 ;
        RECT  5.170 1.025 5.330 1.555 ;
        RECT  3.730 1.025 5.170 1.185 ;
        RECT  3.470 1.025 3.730 1.535 ;
        RECT  2.030 1.025 3.470 1.185 ;
        RECT  1.770 1.025 2.030 1.540 ;
        RECT  0.335 1.025 1.770 1.185 ;
        RECT  0.160 1.025 0.335 2.400 ;
        RECT  0.125 1.515 0.160 2.400 ;
        END
        ANTENNAGATEAREA     1.4976 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.200 -0.250 12.880 0.250 ;
        RECT  11.940 -0.250 12.200 0.405 ;
        RECT  10.500 -0.250 11.940 0.250 ;
        RECT  10.240 -0.250 10.500 0.405 ;
        RECT  8.605 -0.250 10.240 0.250 ;
        RECT  8.345 -0.250 8.605 0.405 ;
        RECT  6.720 -0.250 8.345 0.250 ;
        RECT  6.460 -0.250 6.720 0.405 ;
        RECT  5.630 -0.250 6.460 0.250 ;
        RECT  5.370 -0.250 5.630 0.405 ;
        RECT  3.930 -0.250 5.370 0.250 ;
        RECT  3.670 -0.250 3.930 0.405 ;
        RECT  2.225 -0.250 3.670 0.250 ;
        RECT  1.965 -0.250 2.225 0.405 ;
        RECT  0.555 -0.250 1.965 0.250 ;
        RECT  0.295 -0.250 0.555 0.755 ;
        RECT  0.000 -0.250 0.295 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.990 3.440 12.880 3.940 ;
        RECT  11.730 3.285 11.990 3.940 ;
        RECT  10.260 3.440 11.730 3.940 ;
        RECT  10.000 3.285 10.260 3.940 ;
        RECT  8.560 3.440 10.000 3.940 ;
        RECT  8.300 3.285 8.560 3.940 ;
        RECT  6.705 3.440 8.300 3.940 ;
        RECT  6.445 3.285 6.705 3.940 ;
        RECT  5.475 3.440 6.445 3.940 ;
        RECT  5.215 3.285 5.475 3.940 ;
        RECT  3.760 3.440 5.215 3.940 ;
        RECT  3.500 3.285 3.760 3.940 ;
        RECT  2.060 3.440 3.500 3.940 ;
        RECT  1.800 3.285 2.060 3.940 ;
        RECT  0.385 3.440 1.800 3.940 ;
        RECT  0.335 2.935 0.385 3.940 ;
        RECT  0.125 2.595 0.335 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.930 1.755 11.030 1.915 ;
        RECT  10.770 1.755 10.930 2.585 ;
        RECT  9.340 2.425 10.770 2.585 ;
        RECT  9.080 1.755 9.340 2.585 ;
        RECT  7.880 2.425 9.080 2.585 ;
        RECT  7.620 1.705 7.880 2.585 ;
        RECT  0.675 2.425 7.620 2.585 ;
        RECT  5.770 1.025 6.180 1.185 ;
        RECT  5.610 1.025 5.770 1.895 ;
        RECT  4.940 1.735 5.610 1.895 ;
        RECT  4.780 1.365 4.940 1.895 ;
        RECT  4.680 1.365 4.780 1.645 ;
        RECT  4.070 1.365 4.680 1.525 ;
        RECT  3.910 1.365 4.070 1.875 ;
        RECT  3.245 1.715 3.910 1.875 ;
        RECT  3.085 1.365 3.245 1.875 ;
        RECT  2.985 1.365 3.085 1.595 ;
        RECT  2.370 1.365 2.985 1.525 ;
        RECT  2.210 1.365 2.370 1.900 ;
        RECT  1.495 1.740 2.210 1.900 ;
        RECT  1.335 1.365 1.495 1.900 ;
        RECT  0.675 1.365 1.335 1.525 ;
        RECT  0.515 1.365 0.675 2.585 ;
    END
END MXI2X6

MACRO MXI2X4
    CLASS CORE ;
    FOREIGN MXI2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.065 0.840 5.235 1.135 ;
        RECT  4.975 0.840 5.065 2.215 ;
        RECT  4.855 0.930 4.975 2.215 ;
        RECT  4.210 0.930 4.855 1.135 ;
        RECT  4.805 1.705 4.855 2.215 ;
        RECT  4.045 1.705 4.805 1.905 ;
        RECT  4.140 0.790 4.210 1.135 ;
        RECT  3.950 0.475 4.140 1.135 ;
        RECT  4.015 1.705 4.045 2.740 ;
        RECT  3.785 1.700 4.015 2.740 ;
        RECT  3.190 0.475 3.950 0.665 ;
        RECT  2.765 2.540 3.785 2.740 ;
        RECT  2.930 0.475 3.190 0.795 ;
        END
        ANTENNADIFFAREA     1.9160 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 2.930 5.395 3.220 ;
        RECT  4.910 2.945 5.185 3.220 ;
        RECT  0.925 2.945 4.910 3.105 ;
        RECT  0.665 2.735 0.925 3.105 ;
        END
        ANTENNAGATEAREA     0.7670 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.290 2.175 1.580 ;
        RECT  1.965 1.290 2.150 1.585 ;
        RECT  1.695 1.420 1.965 1.585 ;
        RECT  1.435 1.420 1.695 1.680 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.575 6.435 1.835 ;
        RECT  5.645 1.575 5.855 1.990 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.265 -0.250 6.900 0.250 ;
        RECT  6.005 -0.250 6.265 1.045 ;
        RECT  2.130 -0.250 6.005 0.250 ;
        RECT  1.870 -0.250 2.130 0.405 ;
        RECT  1.325 -0.250 1.870 0.250 ;
        RECT  1.065 -0.250 1.325 0.405 ;
        RECT  0.385 -0.250 1.065 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.265 3.440 6.900 3.940 ;
        RECT  6.005 2.595 6.265 3.940 ;
        RECT  2.285 3.440 6.005 3.940 ;
        RECT  2.025 3.285 2.285 3.940 ;
        RECT  1.185 3.440 2.025 3.940 ;
        RECT  0.925 3.285 1.185 3.940 ;
        RECT  0.385 3.440 0.925 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.615 0.695 6.775 3.195 ;
        RECT  6.515 0.695 6.615 1.395 ;
        RECT  6.515 2.170 6.615 3.195 ;
        RECT  5.750 1.235 6.515 1.395 ;
        RECT  5.755 2.170 6.515 2.330 ;
        RECT  5.495 2.170 5.755 2.750 ;
        RECT  5.650 0.770 5.750 1.395 ;
        RECT  5.590 0.470 5.650 1.395 ;
        RECT  5.490 0.470 5.590 1.030 ;
        RECT  4.555 2.590 5.495 2.750 ;
        RECT  4.720 0.470 5.490 0.630 ;
        RECT  4.460 0.470 4.720 0.745 ;
        RECT  4.295 2.130 4.555 2.750 ;
        RECT  4.290 1.315 4.550 1.520 ;
        RECT  2.805 1.360 4.290 1.520 ;
        RECT  3.440 0.845 3.700 1.165 ;
        RECT  3.275 1.955 3.535 2.360 ;
        RECT  2.680 1.005 3.440 1.165 ;
        RECT  1.735 2.200 3.275 2.360 ;
        RECT  2.645 1.360 2.805 2.020 ;
        RECT  2.420 0.790 2.680 1.165 ;
        RECT  2.500 1.730 2.645 2.020 ;
        RECT  0.785 1.860 2.500 2.020 ;
        RECT  1.725 0.795 2.420 0.955 ;
        RECT  1.475 2.200 1.735 2.750 ;
        RECT  1.625 0.790 1.725 1.050 ;
        RECT  1.465 0.585 1.625 1.050 ;
        RECT  0.260 2.395 1.475 2.555 ;
        RECT  0.260 0.585 1.465 0.745 ;
        RECT  0.625 1.005 0.785 2.215 ;
        RECT  0.525 1.005 0.625 1.265 ;
        RECT  0.525 1.955 0.625 2.215 ;
        RECT  0.100 0.585 0.260 2.555 ;
    END
END MXI2X4

MACRO MXI2X2
    CLASS CORE ;
    FOREIGN MXI2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.355 2.695 3.455 2.955 ;
        RECT  3.195 1.840 3.355 2.955 ;
        RECT  3.005 1.840 3.195 2.000 ;
        RECT  3.095 2.795 3.195 2.955 ;
        RECT  2.885 2.795 3.095 3.220 ;
        RECT  2.845 0.810 3.005 2.000 ;
        RECT  2.430 2.795 2.885 2.955 ;
        RECT  2.745 0.810 2.845 1.070 ;
        RECT  2.270 2.525 2.430 2.955 ;
        RECT  2.170 2.525 2.270 2.785 ;
        END
        ANTENNADIFFAREA     0.8892 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.415 0.795 1.990 ;
        RECT  0.475 1.415 0.585 1.675 ;
        END
        ANTENNAGATEAREA     0.3627 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 1.130 1.715 1.635 ;
        END
        ANTENNAGATEAREA     0.2678 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.305 1.700 4.475 1.990 ;
        RECT  4.145 1.360 4.305 1.990 ;
        RECT  4.045 1.360 4.145 1.620 ;
        END
        ANTENNAGATEAREA     0.2574 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.335 -0.250 4.600 0.250 ;
        RECT  4.075 -0.250 4.335 1.135 ;
        RECT  1.660 -0.250 4.075 0.250 ;
        RECT  0.720 -0.250 1.660 0.795 ;
        RECT  0.000 -0.250 0.720 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 3.440 4.600 3.940 ;
        RECT  4.215 2.200 4.475 3.940 ;
        RECT  1.920 3.440 4.215 3.940 ;
        RECT  1.660 2.520 1.920 3.940 ;
        RECT  0.900 3.440 1.660 3.940 ;
        RECT  0.640 2.295 0.900 3.940 ;
        RECT  0.000 3.440 0.640 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.790 2.275 3.965 3.215 ;
        RECT  3.705 0.575 3.790 3.215 ;
        RECT  3.630 0.575 3.705 2.435 ;
        RECT  3.530 0.575 3.630 1.175 ;
        RECT  3.350 1.355 3.450 1.615 ;
        RECT  3.190 0.470 3.350 1.615 ;
        RECT  2.055 0.470 3.190 0.630 ;
        RECT  2.775 2.355 2.940 2.615 ;
        RECT  2.615 2.180 2.775 2.615 ;
        RECT  2.495 2.180 2.615 2.340 ;
        RECT  2.335 0.810 2.495 2.340 ;
        RECT  2.235 0.810 2.335 1.070 ;
        RECT  1.410 2.180 2.335 2.340 ;
        RECT  2.055 1.740 2.155 2.000 ;
        RECT  1.895 0.470 2.055 2.000 ;
        RECT  1.135 1.840 1.895 2.000 ;
        RECT  1.150 2.180 1.410 2.555 ;
        RECT  0.975 1.075 1.135 2.000 ;
        RECT  0.385 1.075 0.975 1.235 ;
        RECT  0.285 0.975 0.385 1.235 ;
        RECT  0.285 2.205 0.385 2.465 ;
        RECT  0.125 0.975 0.285 2.465 ;
    END
END MXI2X2

MACRO MXI2X1
    CLASS CORE ;
    FOREIGN MXI2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.510 2.635 2.810 ;
        RECT  2.305 2.510 2.425 2.670 ;
        RECT  2.145 0.580 2.305 2.670 ;
        RECT  2.075 0.580 2.145 0.740 ;
        RECT  1.920 2.410 2.145 2.670 ;
        RECT  1.815 0.480 2.075 0.740 ;
        END
        ANTENNADIFFAREA     0.6371 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 2.850 2.245 3.110 ;
        RECT  1.740 2.850 1.985 3.010 ;
        RECT  1.580 2.550 1.740 3.010 ;
        RECT  0.585 2.550 1.580 2.710 ;
        RECT  0.535 2.450 0.585 2.710 ;
        RECT  0.325 2.450 0.535 2.810 ;
        RECT  0.125 2.520 0.325 2.810 ;
        END
        ANTENNAGATEAREA     0.1898 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.935 1.605 1.195 1.865 ;
        RECT  0.795 1.700 0.935 1.865 ;
        RECT  0.585 1.700 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.290 3.095 1.955 ;
        RECT  2.825 1.695 2.885 1.955 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.220 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.955 -0.250 2.835 0.250 ;
        RECT  0.695 -0.250 0.955 1.080 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.220 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.990 3.440 2.835 3.940 ;
        RECT  0.730 2.895 0.990 3.940 ;
        RECT  0.000 3.440 0.730 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.485 0.990 2.645 2.330 ;
        RECT  1.805 0.920 1.965 2.230 ;
        RECT  1.500 0.920 1.805 1.080 ;
        RECT  1.595 2.070 1.805 2.230 ;
        RECT  1.570 1.630 1.625 1.890 ;
        RECT  1.335 2.070 1.595 2.330 ;
        RECT  1.410 1.260 1.570 1.890 ;
        RECT  1.240 0.820 1.500 1.080 ;
        RECT  0.385 1.260 1.410 1.420 ;
        RECT  0.225 0.940 0.385 2.270 ;
        RECT  0.125 0.940 0.225 1.200 ;
        RECT  0.125 2.010 0.225 2.270 ;
    END
END MXI2X1

MACRO MXI2XL
    CLASS CORE ;
    FOREIGN MXI2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.435 2.635 2.810 ;
        RECT  2.265 2.435 2.425 2.595 ;
        RECT  2.105 0.615 2.265 2.595 ;
        RECT  1.835 0.615 2.105 0.775 ;
        RECT  1.800 2.435 2.105 2.595 ;
        RECT  1.540 2.435 1.800 2.785 ;
        END
        ANTENNADIFFAREA     0.4538 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.980 2.865 2.240 3.125 ;
        RECT  1.360 2.965 1.980 3.125 ;
        RECT  1.200 2.495 1.360 3.125 ;
        RECT  0.585 2.495 1.200 2.655 ;
        RECT  0.335 2.395 0.585 2.655 ;
        RECT  0.125 2.395 0.335 2.810 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.635 1.155 1.795 ;
        RECT  0.610 1.635 0.795 1.990 ;
        RECT  0.585 1.700 0.610 1.990 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.080 3.095 1.755 ;
        RECT  2.795 1.495 2.885 1.755 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.220 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.955 -0.250 2.835 0.250 ;
        RECT  0.695 -0.250 0.955 1.115 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.220 3.940 ;
        RECT  2.835 2.895 3.095 3.940 ;
        RECT  0.970 3.440 2.835 3.940 ;
        RECT  0.710 2.895 0.970 3.940 ;
        RECT  0.000 3.440 0.710 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.455 0.995 2.615 2.255 ;
        RECT  1.765 0.955 1.925 2.205 ;
        RECT  1.525 0.955 1.765 1.115 ;
        RECT  1.110 2.045 1.765 2.205 ;
        RECT  1.495 1.585 1.585 1.845 ;
        RECT  1.265 0.855 1.525 1.115 ;
        RECT  1.335 1.295 1.495 1.845 ;
        RECT  0.385 1.295 1.335 1.455 ;
        RECT  0.225 0.855 0.385 2.215 ;
        RECT  0.125 0.855 0.225 1.115 ;
        RECT  0.125 1.955 0.225 2.215 ;
    END
END MXI2XL

MACRO MX4X4
    CLASS CORE ;
    FOREIGN MX4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.580 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.965 0.695 9.995 3.220 ;
        RECT  9.785 0.585 9.965 3.220 ;
        RECT  9.725 0.585 9.785 3.025 ;
        RECT  9.685 0.585 9.725 1.185 ;
        RECT  9.685 2.085 9.725 3.025 ;
        END
        ANTENNADIFFAREA     0.7980 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.105 1.890 9.270 3.090 ;
        RECT  8.965 1.890 9.105 2.150 ;
        RECT  7.695 2.930 9.105 3.090 ;
        RECT  7.485 2.930 7.695 3.220 ;
        RECT  7.235 2.930 7.485 3.190 ;
        END
        ANTENNAGATEAREA     0.3809 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.380 2.965 5.415 3.225 ;
        RECT  5.155 2.930 5.380 3.225 ;
        RECT  1.715 2.930 5.155 3.090 ;
        RECT  4.905 0.495 4.955 0.755 ;
        RECT  4.695 0.495 4.905 0.760 ;
        RECT  3.995 0.585 4.695 0.760 ;
        RECT  3.835 0.585 3.995 1.670 ;
        RECT  2.450 0.585 3.835 0.745 ;
        RECT  3.670 1.510 3.835 1.670 ;
        RECT  2.085 0.485 2.450 0.745 ;
        RECT  1.185 0.585 2.085 0.745 ;
        RECT  1.230 2.930 1.715 3.220 ;
        RECT  1.185 2.930 1.230 3.090 ;
        RECT  1.025 0.585 1.185 3.090 ;
        END
        ANTENNAGATEAREA     0.7566 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.635 3.095 1.990 ;
        RECT  2.595 1.635 2.780 1.795 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.440 0.425 1.855 ;
        RECT  0.125 1.290 0.335 1.855 ;
        END
        ANTENNAGATEAREA     0.2730 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 1.130 4.475 1.675 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.580 6.790 1.840 ;
        RECT  6.565 1.580 6.775 1.990 ;
        RECT  6.370 1.580 6.565 1.840 ;
        END
        ANTENNAGATEAREA     0.2704 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.455 -0.250 10.580 0.250 ;
        RECT  10.195 -0.250 10.455 1.165 ;
        RECT  9.395 -0.250 10.195 0.250 ;
        RECT  9.135 -0.250 9.395 0.405 ;
        RECT  6.860 -0.250 9.135 0.250 ;
        RECT  6.600 -0.250 6.860 0.405 ;
        RECT  4.145 -0.250 6.600 0.250 ;
        RECT  3.885 -0.250 4.145 0.405 ;
        RECT  3.155 -0.250 3.885 0.250 ;
        RECT  2.895 -0.250 3.155 0.405 ;
        RECT  0.385 -0.250 2.895 0.250 ;
        RECT  0.125 -0.250 0.385 1.080 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.455 3.440 10.580 3.940 ;
        RECT  10.195 2.160 10.455 3.940 ;
        RECT  9.405 3.440 10.195 3.940 ;
        RECT  9.145 3.285 9.405 3.940 ;
        RECT  6.895 3.440 9.145 3.940 ;
        RECT  6.635 3.285 6.895 3.940 ;
        RECT  4.060 3.440 6.635 3.940 ;
        RECT  3.800 3.285 4.060 3.940 ;
        RECT  3.035 3.440 3.800 3.940 ;
        RECT  2.775 3.285 3.035 3.940 ;
        RECT  0.385 3.440 2.775 3.940 ;
        RECT  0.125 2.110 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.395 1.395 9.495 1.655 ;
        RECT  9.235 0.635 9.395 1.655 ;
        RECT  8.485 0.635 9.235 0.795 ;
        RECT  8.895 0.990 8.995 1.250 ;
        RECT  8.765 2.480 8.915 2.740 ;
        RECT  8.765 0.990 8.895 1.595 ;
        RECT  8.735 0.990 8.765 2.740 ;
        RECT  8.605 1.435 8.735 2.740 ;
        RECT  6.760 2.580 8.605 2.740 ;
        RECT  8.385 0.635 8.485 1.235 ;
        RECT  8.385 2.095 8.405 2.355 ;
        RECT  8.225 0.635 8.385 2.355 ;
        RECT  8.145 2.095 8.225 2.355 ;
        RECT  7.925 0.585 7.975 1.235 ;
        RECT  7.765 0.585 7.925 2.355 ;
        RECT  7.715 0.585 7.765 1.235 ;
        RECT  7.605 2.095 7.765 2.355 ;
        RECT  5.800 0.585 7.715 0.745 ;
        RECT  7.410 1.315 7.550 1.575 ;
        RECT  7.310 0.940 7.410 1.575 ;
        RECT  7.150 0.940 7.310 2.385 ;
        RECT  7.035 2.125 7.150 2.385 ;
        RECT  6.600 2.580 6.760 3.090 ;
        RECT  5.845 2.930 6.600 3.090 ;
        RECT  6.185 2.145 6.345 2.745 ;
        RECT  6.185 0.955 6.310 1.215 ;
        RECT  6.085 0.955 6.185 2.745 ;
        RECT  6.025 0.955 6.085 2.305 ;
        RECT  5.685 2.550 5.845 3.090 ;
        RECT  5.700 0.530 5.800 1.130 ;
        RECT  5.540 0.530 5.700 2.360 ;
        RECT  1.975 2.550 5.685 2.710 ;
        RECT  5.420 2.100 5.540 2.360 ;
        RECT  5.055 1.105 5.215 2.355 ;
        RECT  5.045 1.105 5.055 1.265 ;
        RECT  4.350 2.195 5.055 2.355 ;
        RECT  4.785 1.005 5.045 1.265 ;
        RECT  4.715 1.535 4.875 2.015 ;
        RECT  3.640 1.855 4.715 2.015 ;
        RECT  3.485 1.025 3.655 1.285 ;
        RECT  3.485 1.855 3.640 2.370 ;
        RECT  3.325 1.025 3.485 2.370 ;
        RECT  2.295 1.275 3.325 1.435 ;
        RECT  1.945 0.925 2.535 1.085 ;
        RECT  2.385 2.110 2.485 2.370 ;
        RECT  2.225 2.015 2.385 2.370 ;
        RECT  2.135 1.275 2.295 1.825 ;
        RECT  1.945 2.015 2.225 2.175 ;
        RECT  1.535 2.450 1.975 2.710 ;
        RECT  1.785 0.925 1.945 2.175 ;
        RECT  1.375 0.925 1.535 2.710 ;
        RECT  1.365 0.925 1.375 1.185 ;
        RECT  0.685 0.560 0.845 3.125 ;
    END
END MX4X4

MACRO MX4X2
    CLASS CORE ;
    FOREIGN MX4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.120 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.835 0.550 9.995 3.195 ;
        RECT  9.785 0.550 9.835 0.945 ;
        RECT  9.735 2.255 9.835 3.195 ;
        RECT  9.735 0.550 9.785 0.810 ;
        END
        ANTENNADIFFAREA     0.7140 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.490 2.335 9.535 2.810 ;
        RECT  9.485 1.865 9.490 2.810 ;
        RECT  9.325 1.865 9.485 3.095 ;
        RECT  9.125 1.865 9.325 2.025 ;
        RECT  7.555 2.935 9.325 3.095 ;
        RECT  8.965 1.415 9.125 2.025 ;
        RECT  7.295 2.935 7.555 3.195 ;
        END
        ANTENNAGATEAREA     0.3809 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.130 2.930 5.390 3.225 ;
        RECT  1.715 2.930 5.130 3.090 ;
        RECT  4.755 0.495 5.015 0.755 ;
        RECT  3.985 0.585 4.755 0.745 ;
        RECT  3.725 0.585 3.985 0.830 ;
        RECT  3.555 0.585 3.725 0.760 ;
        RECT  2.450 0.585 3.555 0.745 ;
        RECT  2.090 0.485 2.450 0.745 ;
        RECT  1.185 0.535 2.090 0.695 ;
        RECT  1.185 2.930 1.715 3.220 ;
        RECT  1.025 0.535 1.185 3.220 ;
        END
        ANTENNAGATEAREA     0.7566 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.750 1.635 3.095 1.990 ;
        RECT  2.565 1.635 2.750 1.795 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.495 0.455 1.755 ;
        RECT  0.125 1.290 0.335 1.755 ;
        END
        ANTENNAGATEAREA     0.2730 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 1.290 4.475 1.580 ;
        RECT  4.140 1.150 4.440 1.625 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 1.290 6.880 1.840 ;
        RECT  6.400 1.580 6.565 1.840 ;
        END
        ANTENNAGATEAREA     0.2704 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.455 -0.250 10.120 0.250 ;
        RECT  9.195 -0.250 9.455 0.405 ;
        RECT  6.870 -0.250 9.195 0.250 ;
        RECT  6.610 -0.250 6.870 0.405 ;
        RECT  4.205 -0.250 6.610 0.250 ;
        RECT  3.945 -0.250 4.205 0.405 ;
        RECT  3.165 -0.250 3.945 0.250 ;
        RECT  2.905 -0.250 3.165 0.405 ;
        RECT  0.385 -0.250 2.905 0.250 ;
        RECT  0.125 -0.250 0.385 1.080 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.455 3.440 10.120 3.940 ;
        RECT  9.195 3.285 9.455 3.940 ;
        RECT  6.955 3.440 9.195 3.940 ;
        RECT  6.695 3.285 6.955 3.940 ;
        RECT  4.065 3.440 6.695 3.940 ;
        RECT  3.805 3.285 4.065 3.940 ;
        RECT  3.035 3.440 3.805 3.940 ;
        RECT  2.775 3.285 3.035 3.940 ;
        RECT  0.385 3.440 2.775 3.940 ;
        RECT  0.125 2.110 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.555 1.385 9.655 1.645 ;
        RECT  9.395 0.635 9.555 1.645 ;
        RECT  8.545 0.635 9.395 0.795 ;
        RECT  8.795 0.975 9.055 1.235 ;
        RECT  8.775 2.480 8.945 2.740 ;
        RECT  8.775 1.075 8.795 1.235 ;
        RECT  8.615 1.075 8.775 2.740 ;
        RECT  6.790 2.580 8.615 2.740 ;
        RECT  8.435 0.535 8.545 0.795 ;
        RECT  8.275 0.535 8.435 2.355 ;
        RECT  8.175 2.095 8.275 2.355 ;
        RECT  7.925 0.585 8.035 1.200 ;
        RECT  7.765 0.585 7.925 2.355 ;
        RECT  5.810 0.585 7.765 0.745 ;
        RECT  7.665 2.095 7.765 2.355 ;
        RECT  7.420 1.315 7.570 1.575 ;
        RECT  7.355 0.940 7.420 1.575 ;
        RECT  7.195 0.940 7.355 2.385 ;
        RECT  7.160 0.940 7.195 1.540 ;
        RECT  7.095 2.125 7.195 2.385 ;
        RECT  6.630 2.580 6.790 3.090 ;
        RECT  5.770 2.930 6.630 3.090 ;
        RECT  6.220 2.145 6.405 2.745 ;
        RECT  6.220 0.955 6.320 1.215 ;
        RECT  6.145 0.955 6.220 2.745 ;
        RECT  6.060 0.955 6.145 2.395 ;
        RECT  5.710 0.530 5.810 1.130 ;
        RECT  5.610 2.550 5.770 3.090 ;
        RECT  5.710 2.070 5.720 2.330 ;
        RECT  5.550 0.530 5.710 2.330 ;
        RECT  1.975 2.550 5.610 2.710 ;
        RECT  5.460 2.070 5.550 2.330 ;
        RECT  5.250 0.935 5.275 1.195 ;
        RECT  5.090 0.935 5.250 2.355 ;
        RECT  4.675 0.935 5.090 1.195 ;
        RECT  4.355 2.195 5.090 2.355 ;
        RECT  4.745 1.535 4.905 2.015 ;
        RECT  3.620 1.855 4.745 2.015 ;
        RECT  3.620 1.025 3.715 1.285 ;
        RECT  3.460 1.025 3.620 2.215 ;
        RECT  3.455 1.025 3.460 1.435 ;
        RECT  3.325 1.955 3.460 2.215 ;
        RECT  2.285 1.275 3.455 1.435 ;
        RECT  1.920 0.925 2.530 1.085 ;
        RECT  2.225 2.015 2.485 2.275 ;
        RECT  2.125 1.275 2.285 1.690 ;
        RECT  1.920 2.015 2.225 2.175 ;
        RECT  1.530 2.450 1.975 2.710 ;
        RECT  1.760 0.925 1.920 2.175 ;
        RECT  1.370 0.985 1.530 2.710 ;
        RECT  0.685 0.560 0.845 3.125 ;
    END
END MX4X2

MACRO MX4X1
    CLASS CORE ;
    FOREIGN MX4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.600 0.975 8.615 2.810 ;
        RECT  8.440 0.975 8.600 2.935 ;
        RECT  8.430 0.975 8.440 1.355 ;
        RECT  8.340 2.335 8.440 2.935 ;
        RECT  8.355 0.975 8.430 1.235 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 0.510 6.490 0.760 ;
        RECT  6.105 0.470 6.315 0.760 ;
        RECT  5.860 0.510 6.105 0.760 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.530 2.780 1.790 ;
        RECT  2.520 1.290 2.635 1.790 ;
        RECT  2.450 1.290 2.520 1.725 ;
        RECT  2.425 1.290 2.450 1.580 ;
        END
        ANTENNAGATEAREA     0.4472 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 1.255 2.225 1.760 ;
        RECT  1.965 1.290 1.975 1.580 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.635 0.435 1.895 ;
        RECT  0.175 1.290 0.335 1.895 ;
        RECT  0.125 1.290 0.175 1.765 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.070 3.590 1.640 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.645 1.700 5.855 1.990 ;
        RECT  5.385 1.700 5.645 1.860 ;
        RECT  5.225 1.465 5.385 1.860 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.215 -0.250 8.740 0.250 ;
        RECT  7.955 -0.250 8.215 0.405 ;
        RECT  5.600 -0.250 7.955 0.250 ;
        RECT  5.340 -0.250 5.600 0.925 ;
        RECT  3.480 -0.250 5.340 0.250 ;
        RECT  3.220 -0.250 3.480 0.775 ;
        RECT  2.500 -0.250 3.220 0.250 ;
        RECT  2.240 -0.250 2.500 1.070 ;
        RECT  0.385 -0.250 2.240 0.250 ;
        RECT  0.125 -0.250 0.385 1.000 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 3.440 8.740 3.940 ;
        RECT  7.800 3.285 8.060 3.940 ;
        RECT  5.680 3.440 7.800 3.940 ;
        RECT  5.420 3.285 5.680 3.940 ;
        RECT  3.380 3.440 5.420 3.940 ;
        RECT  3.120 3.095 3.380 3.940 ;
        RECT  2.535 3.440 3.120 3.940 ;
        RECT  2.275 3.095 2.535 3.940 ;
        RECT  0.425 3.440 2.275 3.940 ;
        RECT  0.165 3.285 0.425 3.940 ;
        RECT  0.000 3.440 0.165 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.155 1.635 8.255 1.895 ;
        RECT  7.995 0.600 8.155 1.895 ;
        RECT  7.195 0.600 7.995 0.760 ;
        RECT  7.540 0.945 7.705 1.205 ;
        RECT  7.540 2.165 7.640 2.865 ;
        RECT  7.380 0.945 7.540 3.100 ;
        RECT  3.960 2.940 7.380 3.100 ;
        RECT  7.035 0.600 7.195 1.110 ;
        RECT  7.030 2.155 7.130 2.755 ;
        RECT  7.030 0.850 7.035 1.110 ;
        RECT  6.870 0.850 7.030 2.755 ;
        RECT  6.570 0.945 6.685 2.305 ;
        RECT  6.525 0.945 6.570 2.755 ;
        RECT  6.425 0.945 6.525 1.205 ;
        RECT  6.410 2.145 6.525 2.755 ;
        RECT  4.705 2.580 6.410 2.740 ;
        RECT  6.225 1.465 6.330 1.725 ;
        RECT  6.065 0.940 6.225 2.360 ;
        RECT  5.915 0.940 6.065 1.200 ;
        RECT  5.845 2.200 6.065 2.360 ;
        RECT  5.045 0.750 5.050 0.910 ;
        RECT  4.885 0.750 5.045 2.370 ;
        RECT  4.790 0.750 4.885 0.910 ;
        RECT  4.545 1.095 4.705 2.740 ;
        RECT  4.540 1.095 4.545 1.255 ;
        RECT  4.260 2.580 4.545 2.740 ;
        RECT  4.380 0.735 4.540 1.255 ;
        RECT  4.280 0.735 4.380 0.995 ;
        RECT  4.205 1.435 4.365 2.380 ;
        RECT  4.030 1.435 4.205 1.595 ;
        RECT  3.930 2.220 4.205 2.380 ;
        RECT  3.870 0.790 4.030 1.595 ;
        RECT  3.865 1.775 4.025 2.035 ;
        RECT  3.800 2.750 3.960 3.100 ;
        RECT  3.670 2.220 3.930 2.480 ;
        RECT  3.770 0.790 3.870 1.050 ;
        RECT  3.140 1.860 3.865 2.035 ;
        RECT  1.440 2.750 3.800 2.910 ;
        RECT  3.015 1.080 3.140 2.345 ;
        RECT  3.000 1.080 3.015 2.555 ;
        RECT  2.980 1.030 3.000 2.555 ;
        RECT  2.840 1.030 2.980 1.290 ;
        RECT  2.755 2.185 2.980 2.555 ;
        RECT  2.355 2.185 2.755 2.345 ;
        RECT  2.195 1.940 2.355 2.345 ;
        RECT  1.795 1.940 2.195 2.100 ;
        RECT  1.780 0.750 1.990 1.010 ;
        RECT  1.730 2.280 1.990 2.540 ;
        RECT  1.635 1.800 1.795 2.100 ;
        RECT  1.620 0.750 1.780 1.620 ;
        RECT  1.455 2.280 1.730 2.440 ;
        RECT  1.455 1.460 1.620 1.620 ;
        RECT  1.295 1.460 1.455 2.440 ;
        RECT  1.340 0.845 1.440 1.105 ;
        RECT  1.180 2.625 1.440 2.910 ;
        RECT  1.180 0.845 1.340 1.270 ;
        RECT  1.115 1.110 1.180 1.270 ;
        RECT  1.115 2.625 1.180 2.785 ;
        RECT  0.955 1.110 1.115 2.785 ;
        RECT  0.775 0.760 0.930 0.920 ;
        RECT  0.615 0.760 0.775 2.780 ;
    END
END MX4X1

MACRO MX4XL
    CLASS CORE ;
    FOREIGN MX4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.450 0.975 8.615 2.915 ;
        RECT  8.430 0.975 8.450 1.355 ;
        RECT  8.405 2.110 8.450 2.915 ;
        RECT  8.355 0.975 8.430 1.235 ;
        RECT  8.350 2.655 8.405 2.915 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 0.510 6.490 0.760 ;
        RECT  6.105 0.470 6.315 0.760 ;
        RECT  5.860 0.510 6.105 0.760 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.475 2.790 2.050 ;
        RECT  2.630 1.290 2.635 2.050 ;
        RECT  2.425 1.290 2.630 1.635 ;
        END
        ANTENNAGATEAREA     0.1560 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 1.260 2.225 1.750 ;
        RECT  1.965 1.290 1.985 1.580 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.395 1.895 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.000 3.565 1.570 ;
        RECT  3.345 1.000 3.555 1.580 ;
        RECT  3.320 1.000 3.345 1.570 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.830 1.700 5.855 1.990 ;
        RECT  5.645 1.570 5.830 1.990 ;
        RECT  5.490 1.570 5.645 1.730 ;
        RECT  5.230 1.355 5.490 1.730 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.185 -0.250 8.740 0.250 ;
        RECT  7.925 -0.250 8.185 0.405 ;
        RECT  5.620 -0.250 7.925 0.250 ;
        RECT  5.360 -0.250 5.620 0.405 ;
        RECT  3.470 -0.250 5.360 0.250 ;
        RECT  3.210 -0.250 3.470 0.775 ;
        RECT  2.530 -0.250 3.210 0.250 ;
        RECT  2.270 -0.250 2.530 1.075 ;
        RECT  0.385 -0.250 2.270 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.100 3.440 8.740 3.940 ;
        RECT  7.840 2.645 8.100 3.940 ;
        RECT  7.810 3.285 7.840 3.940 ;
        RECT  5.665 3.440 7.810 3.940 ;
        RECT  5.405 3.285 5.665 3.940 ;
        RECT  3.360 3.440 5.405 3.940 ;
        RECT  3.100 3.095 3.360 3.940 ;
        RECT  2.420 3.440 3.100 3.940 ;
        RECT  2.160 3.095 2.420 3.940 ;
        RECT  0.385 3.440 2.160 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.175 1.635 8.270 1.895 ;
        RECT  8.015 0.660 8.175 1.895 ;
        RECT  7.245 0.660 8.015 0.820 ;
        RECT  8.010 1.635 8.015 1.895 ;
        RECT  7.655 2.135 7.755 2.395 ;
        RECT  7.655 1.025 7.675 1.285 ;
        RECT  7.495 1.025 7.655 3.030 ;
        RECT  7.415 1.025 7.495 1.285 ;
        RECT  4.060 2.870 7.495 3.030 ;
        RECT  7.185 0.560 7.245 0.820 ;
        RECT  7.025 0.560 7.185 2.395 ;
        RECT  6.985 0.560 7.025 0.820 ;
        RECT  6.925 2.135 7.025 2.395 ;
        RECT  6.600 1.010 6.710 1.270 ;
        RECT  6.440 1.010 6.600 2.690 ;
        RECT  6.405 2.135 6.440 2.690 ;
        RECT  4.695 2.530 6.405 2.690 ;
        RECT  6.225 1.410 6.260 1.670 ;
        RECT  6.065 0.940 6.225 2.350 ;
        RECT  5.940 0.940 6.065 1.200 ;
        RECT  5.845 2.190 6.065 2.350 ;
        RECT  5.035 0.905 5.190 1.165 ;
        RECT  4.875 0.905 5.035 2.315 ;
        RECT  4.535 0.845 4.695 2.690 ;
        RECT  4.360 0.845 4.535 1.105 ;
        RECT  4.250 2.445 4.535 2.690 ;
        RECT  4.195 1.285 4.355 2.265 ;
        RECT  4.050 1.285 4.195 1.445 ;
        RECT  3.940 2.105 4.195 2.265 ;
        RECT  3.900 2.725 4.060 3.030 ;
        RECT  3.890 0.905 4.050 1.445 ;
        RECT  3.855 1.625 4.015 1.925 ;
        RECT  3.680 2.105 3.940 2.405 ;
        RECT  1.385 2.725 3.900 2.885 ;
        RECT  3.790 0.905 3.890 1.165 ;
        RECT  3.130 1.760 3.855 1.925 ;
        RECT  3.000 1.030 3.130 2.440 ;
        RECT  2.970 1.030 3.000 2.490 ;
        RECT  2.840 1.030 2.970 1.290 ;
        RECT  2.740 2.230 2.970 2.490 ;
        RECT  2.315 2.230 2.740 2.390 ;
        RECT  2.155 1.935 2.315 2.390 ;
        RECT  1.795 1.935 2.155 2.095 ;
        RECT  1.785 0.820 1.960 1.080 ;
        RECT  1.695 2.280 1.955 2.540 ;
        RECT  1.635 1.815 1.795 2.095 ;
        RECT  1.700 0.820 1.785 1.630 ;
        RECT  1.625 0.920 1.700 1.630 ;
        RECT  1.455 2.280 1.695 2.440 ;
        RECT  1.455 1.470 1.625 1.630 ;
        RECT  1.295 1.470 1.455 2.440 ;
        RECT  1.130 1.030 1.390 1.290 ;
        RECT  1.115 2.620 1.385 2.885 ;
        RECT  1.115 1.130 1.130 1.290 ;
        RECT  0.955 1.130 1.115 2.885 ;
        RECT  0.605 1.030 0.765 2.445 ;
    END
END MX4XL

MACRO MX2X8
    CLASS CORE ;
    FOREIGN MX2X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.345 0.695 5.395 2.995 ;
        RECT  5.085 0.580 5.345 3.120 ;
        RECT  4.725 0.920 5.085 2.400 ;
        RECT  4.325 0.920 4.725 1.330 ;
        RECT  4.275 2.000 4.725 2.400 ;
        RECT  4.065 0.580 4.325 1.330 ;
        RECT  4.115 2.000 4.275 3.120 ;
        END
        ANTENNADIFFAREA     1.6112 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.305 3.055 1.635 3.215 ;
        RECT  1.145 2.490 1.305 3.215 ;
        RECT  1.045 2.490 1.145 2.995 ;
        RECT  0.395 2.490 1.045 2.650 ;
        RECT  0.335 2.490 0.395 2.795 ;
        RECT  0.125 2.490 0.335 2.810 ;
        END
        ANTENNAGATEAREA     0.3809 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.990 0.880 1.255 1.480 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.255 3.595 2.075 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 -0.250 5.980 0.250 ;
        RECT  5.595 -0.250 5.855 1.075 ;
        RECT  4.835 -0.250 5.595 0.250 ;
        RECT  4.575 -0.250 4.835 0.735 ;
        RECT  3.815 -0.250 4.575 0.250 ;
        RECT  3.555 -0.250 3.815 1.075 ;
        RECT  1.285 -0.250 3.555 0.250 ;
        RECT  1.025 -0.250 1.285 0.700 ;
        RECT  0.000 -0.250 1.025 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 3.440 5.980 3.940 ;
        RECT  5.595 2.255 5.855 3.940 ;
        RECT  4.835 3.440 5.595 3.940 ;
        RECT  4.575 2.595 4.835 3.940 ;
        RECT  3.815 3.440 4.575 3.940 ;
        RECT  3.555 2.935 3.815 3.940 ;
        RECT  0.835 3.440 3.555 3.940 ;
        RECT  0.575 2.880 0.835 3.940 ;
        RECT  0.000 3.440 0.575 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.945 1.560 4.205 1.820 ;
        RECT  3.935 1.660 3.945 1.820 ;
        RECT  3.775 1.660 3.935 2.755 ;
        RECT  2.795 2.595 3.775 2.755 ;
        RECT  3.165 0.475 3.305 1.075 ;
        RECT  3.165 2.255 3.305 2.415 ;
        RECT  3.045 0.475 3.165 2.415 ;
        RECT  3.005 0.915 3.045 2.415 ;
        RECT  2.665 0.550 2.825 1.585 ;
        RECT  2.745 2.485 2.795 2.755 ;
        RECT  2.695 2.485 2.745 2.875 ;
        RECT  2.535 1.790 2.695 2.875 ;
        RECT  1.630 0.550 2.665 0.710 ;
        RECT  2.485 1.790 2.535 1.950 ;
        RECT  1.845 2.715 2.535 2.875 ;
        RECT  2.325 0.930 2.485 1.950 ;
        RECT  2.145 2.150 2.285 2.535 ;
        RECT  2.025 0.995 2.145 2.535 ;
        RECT  1.985 0.995 2.025 2.310 ;
        RECT  1.970 0.995 1.985 1.155 ;
        RECT  1.375 2.150 1.985 2.310 ;
        RECT  1.810 0.895 1.970 1.155 ;
        RECT  1.685 2.535 1.845 2.875 ;
        RECT  1.645 1.660 1.805 1.970 ;
        RECT  1.515 2.535 1.685 2.695 ;
        RECT  1.630 1.660 1.645 1.820 ;
        RECT  1.470 0.550 1.630 1.820 ;
        RECT  0.405 1.660 1.470 1.820 ;
        RECT  1.115 2.005 1.375 2.310 ;
        RECT  0.480 0.580 0.740 0.840 ;
        RECT  0.405 0.650 0.480 0.840 ;
        RECT  0.245 0.650 0.405 2.215 ;
        RECT  0.145 1.955 0.245 2.215 ;
    END
END MX2X8

MACRO MX2X6
    CLASS CORE ;
    FOREIGN MX2X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.390 0.695 5.395 2.995 ;
        RECT  5.130 0.675 5.390 3.120 ;
        RECT  4.725 1.095 5.130 2.400 ;
        RECT  4.370 1.095 4.725 1.395 ;
        RECT  4.370 2.100 4.725 2.400 ;
        RECT  4.110 0.675 4.370 1.395 ;
        RECT  4.110 2.100 4.370 3.045 ;
        END
        ANTENNADIFFAREA     1.5264 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.440 3.000 1.600 3.260 ;
        RECT  1.350 3.000 1.440 3.160 ;
        RECT  1.190 2.520 1.350 3.160 ;
        RECT  0.440 2.520 1.190 2.680 ;
        RECT  0.125 2.520 0.440 2.810 ;
        END
        ANTENNAGATEAREA     0.3809 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.455 1.270 1.615 ;
        RECT  0.610 1.290 0.795 1.615 ;
        RECT  0.585 1.290 0.610 1.580 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.255 3.590 2.075 ;
        END
        ANTENNAGATEAREA     0.2782 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 -0.250 5.520 0.250 ;
        RECT  4.620 -0.250 4.880 0.735 ;
        RECT  3.860 -0.250 4.620 0.250 ;
        RECT  3.600 -0.250 3.860 1.075 ;
        RECT  1.295 -0.250 3.600 0.250 ;
        RECT  1.035 -0.250 1.295 0.930 ;
        RECT  0.000 -0.250 1.035 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 3.440 5.520 3.940 ;
        RECT  4.620 2.595 4.880 3.940 ;
        RECT  3.860 3.440 4.620 3.940 ;
        RECT  3.600 2.935 3.860 3.940 ;
        RECT  0.880 3.440 3.600 3.940 ;
        RECT  0.620 2.880 0.880 3.940 ;
        RECT  0.000 3.440 0.620 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.990 1.575 4.250 1.835 ;
        RECT  3.930 1.675 3.990 1.835 ;
        RECT  3.770 1.675 3.930 2.755 ;
        RECT  2.790 2.595 3.770 2.755 ;
        RECT  3.165 0.475 3.350 1.075 ;
        RECT  3.165 2.255 3.350 2.415 ;
        RECT  3.090 0.475 3.165 2.415 ;
        RECT  3.005 0.915 3.090 2.415 ;
        RECT  2.665 0.550 2.825 1.535 ;
        RECT  2.630 1.790 2.790 2.925 ;
        RECT  1.635 0.550 2.665 0.710 ;
        RECT  2.560 1.375 2.665 1.535 ;
        RECT  2.380 1.790 2.630 1.950 ;
        RECT  1.940 2.765 2.630 2.925 ;
        RECT  2.380 0.930 2.485 1.190 ;
        RECT  2.220 0.930 2.380 1.950 ;
        RECT  2.120 2.135 2.280 2.585 ;
        RECT  2.040 2.135 2.120 2.310 ;
        RECT  1.880 0.895 2.040 2.310 ;
        RECT  1.780 2.660 1.940 2.925 ;
        RECT  1.815 0.895 1.880 1.155 ;
        RECT  1.160 2.150 1.880 2.310 ;
        RECT  1.530 2.660 1.780 2.820 ;
        RECT  1.635 1.710 1.700 1.970 ;
        RECT  1.475 0.550 1.635 1.970 ;
        RECT  0.385 1.810 1.475 1.970 ;
        RECT  0.525 0.700 0.785 0.960 ;
        RECT  0.385 0.800 0.525 0.960 ;
        RECT  0.225 0.800 0.385 2.215 ;
        RECT  0.125 1.955 0.225 2.215 ;
    END
END MX2X6

MACRO MX2X4
    CLASS CORE ;
    FOREIGN MX2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.840 0.880 4.935 1.580 ;
        RECT  4.780 2.115 4.885 2.375 ;
        RECT  4.780 0.675 4.840 1.580 ;
        RECT  4.580 0.675 4.780 2.375 ;
        END
        ANTENNADIFFAREA     0.7642 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.735 0.445 2.995 ;
        RECT  0.125 2.520 0.335 2.995 ;
        END
        ANTENNAGATEAREA     0.3705 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.625 1.065 1.990 ;
        END
        ANTENNAGATEAREA     0.2808 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.980 1.290 4.015 1.580 ;
        RECT  3.805 1.290 3.980 1.895 ;
        RECT  3.730 1.445 3.805 1.895 ;
        END
        ANTENNAGATEAREA     0.2626 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.385 -0.250 5.520 0.250 ;
        RECT  5.125 -0.250 5.385 1.180 ;
        RECT  4.300 -0.250 5.125 0.250 ;
        RECT  4.040 -0.250 4.300 0.755 ;
        RECT  0.925 -0.250 4.040 0.250 ;
        RECT  0.665 -0.250 0.925 1.075 ;
        RECT  0.000 -0.250 0.665 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 3.440 5.520 3.940 ;
        RECT  5.135 2.910 5.395 3.940 ;
        RECT  4.375 3.440 5.135 3.940 ;
        RECT  4.115 2.910 4.375 3.940 ;
        RECT  1.935 3.440 4.115 3.940 ;
        RECT  1.675 2.220 1.935 3.940 ;
        RECT  0.915 3.440 1.675 3.940 ;
        RECT  0.655 2.200 0.915 3.940 ;
        RECT  0.000 3.440 0.655 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.095 1.770 5.255 2.715 ;
        RECT  4.975 1.770 5.095 1.930 ;
        RECT  3.355 2.555 5.095 2.715 ;
        RECT  4.210 0.950 4.370 2.255 ;
        RECT  3.710 0.950 4.210 1.110 ;
        RECT  3.865 2.095 4.210 2.255 ;
        RECT  3.605 2.095 3.865 2.355 ;
        RECT  3.550 0.775 3.710 1.110 ;
        RECT  3.210 0.470 3.370 1.665 ;
        RECT  3.240 2.405 3.355 3.005 ;
        RECT  3.080 1.960 3.240 3.185 ;
        RECT  1.265 0.470 3.210 0.630 ;
        RECT  3.030 1.960 3.080 2.120 ;
        RECT  2.285 3.025 3.080 3.185 ;
        RECT  2.870 0.930 3.030 2.120 ;
        RECT  2.745 2.585 2.845 2.845 ;
        RECT  2.585 2.370 2.745 2.845 ;
        RECT  2.400 2.370 2.585 2.535 ;
        RECT  2.400 0.850 2.570 1.110 ;
        RECT  2.310 0.850 2.400 2.535 ;
        RECT  2.240 0.935 2.310 2.535 ;
        RECT  2.125 2.745 2.285 3.185 ;
        RECT  1.705 0.935 2.240 1.095 ;
        RECT  1.425 1.875 2.240 2.035 ;
        RECT  1.745 1.285 2.005 1.670 ;
        RECT  1.265 1.285 1.745 1.445 ;
        RECT  1.445 0.835 1.705 1.095 ;
        RECT  1.265 1.875 1.425 2.770 ;
        RECT  1.105 0.470 1.265 1.445 ;
        RECT  1.165 2.170 1.265 2.770 ;
        RECT  0.395 1.285 1.105 1.445 ;
        RECT  0.385 1.035 0.395 1.445 ;
        RECT  0.225 1.035 0.385 2.310 ;
        RECT  0.125 1.035 0.225 1.295 ;
        RECT  0.125 2.050 0.225 2.310 ;
    END
END MX2X4

MACRO MX2X2
    CLASS CORE ;
    FOREIGN MX2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 1.290 4.015 2.585 ;
        RECT  3.805 1.130 3.970 3.010 ;
        RECT  3.545 0.695 3.805 1.295 ;
        RECT  3.695 1.990 3.805 3.010 ;
        END
        ANTENNADIFFAREA     0.7460 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 2.705 0.515 2.965 ;
        RECT  0.125 2.705 0.420 3.220 ;
        END
        ANTENNAGATEAREA     0.2951 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.705 1.155 1.925 ;
        RECT  0.585 1.700 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.825 1.155 3.095 1.665 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 -0.250 4.140 0.250 ;
        RECT  2.975 -0.250 3.235 0.875 ;
        RECT  0.985 -0.250 2.975 0.250 ;
        RECT  0.725 -0.250 0.985 0.950 ;
        RECT  0.000 -0.250 0.725 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.415 3.440 4.140 3.940 ;
        RECT  3.155 2.215 3.415 3.940 ;
        RECT  0.955 3.440 3.155 3.940 ;
        RECT  0.695 2.405 0.955 3.940 ;
        RECT  0.000 3.440 0.695 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.515 1.510 3.625 1.770 ;
        RECT  3.355 1.510 3.515 2.035 ;
        RECT  2.975 1.875 3.355 2.035 ;
        RECT  2.815 1.875 2.975 2.895 ;
        RECT  2.265 2.735 2.815 2.895 ;
        RECT  2.475 0.690 2.635 2.555 ;
        RECT  2.105 0.680 2.265 2.895 ;
        RECT  1.835 0.680 2.105 0.840 ;
        RECT  1.845 2.480 2.105 2.740 ;
        RECT  1.765 1.020 1.925 2.300 ;
        RECT  1.525 1.020 1.765 1.180 ;
        RECT  1.525 2.140 1.765 2.300 ;
        RECT  1.425 1.360 1.585 1.930 ;
        RECT  1.265 0.920 1.525 1.180 ;
        RECT  1.265 2.140 1.525 2.835 ;
        RECT  0.405 1.360 1.425 1.520 ;
        RECT  0.405 2.170 0.415 2.430 ;
        RECT  0.245 1.035 0.405 2.430 ;
        RECT  0.125 1.035 0.245 1.295 ;
        RECT  0.155 2.170 0.245 2.430 ;
    END
END MX2X2

MACRO MX2X1
    CLASS CORE ;
    FOREIGN MX2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 0.870 3.555 2.810 ;
        RECT  3.345 0.870 3.395 1.355 ;
        RECT  3.370 2.335 3.395 2.810 ;
        RECT  3.345 2.350 3.370 2.810 ;
        RECT  3.295 0.870 3.345 1.130 ;
        RECT  3.295 2.350 3.345 2.800 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.435 2.725 0.485 2.985 ;
        RECT  0.335 2.725 0.435 3.210 ;
        RECT  0.225 2.725 0.335 3.220 ;
        RECT  0.125 2.930 0.225 3.220 ;
        END
        ANTENNAGATEAREA     0.1560 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.960 1.065 2.220 ;
        RECT  0.585 1.960 0.795 2.400 ;
        RECT  0.580 1.960 0.585 2.220 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.695 1.170 3.095 1.580 ;
        END
        ANTENNAGATEAREA     0.1066 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 -0.250 3.680 0.250 ;
        RECT  2.865 -0.250 3.125 0.405 ;
        RECT  0.955 -0.250 2.865 0.250 ;
        RECT  0.695 -0.250 0.955 1.065 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.150 3.440 3.680 3.940 ;
        RECT  2.890 3.285 3.150 3.940 ;
        RECT  0.955 3.440 2.890 3.940 ;
        RECT  0.695 2.585 0.955 3.940 ;
        RECT  0.000 3.440 0.695 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.080 1.785 3.200 2.045 ;
        RECT  2.920 1.785 3.080 2.935 ;
        RECT  2.175 2.775 2.920 2.935 ;
        RECT  2.355 0.785 2.515 2.595 ;
        RECT  2.015 0.835 2.175 2.935 ;
        RECT  1.715 0.835 2.015 0.995 ;
        RECT  1.715 2.440 2.015 2.700 ;
        RECT  1.675 1.185 1.835 2.260 ;
        RECT  1.465 1.185 1.675 1.345 ;
        RECT  1.465 2.100 1.675 2.260 ;
        RECT  1.335 1.535 1.495 1.795 ;
        RECT  1.305 0.805 1.465 1.345 ;
        RECT  1.305 2.100 1.465 2.660 ;
        RECT  0.385 1.535 1.335 1.695 ;
        RECT  1.205 0.805 1.305 1.065 ;
        RECT  1.205 2.400 1.305 2.660 ;
        RECT  0.225 0.875 0.385 2.520 ;
        RECT  0.125 0.875 0.225 1.135 ;
        RECT  0.125 2.260 0.225 2.520 ;
    END
END MX2X1

MACRO MX2XL
    CLASS CORE ;
    FOREIGN MX2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 0.885 3.565 2.745 ;
        RECT  3.405 0.885 3.555 2.810 ;
        RECT  3.345 0.885 3.405 1.355 ;
        RECT  3.370 2.335 3.405 2.810 ;
        RECT  3.345 2.345 3.370 2.810 ;
        RECT  3.295 0.885 3.345 1.145 ;
        RECT  3.295 2.345 3.345 2.795 ;
        END
        ANTENNADIFFAREA     0.2330 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.725 0.485 3.210 ;
        RECT  0.225 2.725 0.335 3.220 ;
        RECT  0.125 2.930 0.225 3.220 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 2.015 1.125 2.275 ;
        RECT  0.585 2.015 0.795 2.400 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.665 1.170 3.095 1.580 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 -0.250 3.680 0.250 ;
        RECT  2.865 -0.250 3.125 0.405 ;
        RECT  0.955 -0.250 2.865 0.250 ;
        RECT  0.695 -0.250 0.955 1.065 ;
        RECT  0.000 -0.250 0.695 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 3.440 3.680 3.940 ;
        RECT  2.895 3.285 3.155 3.940 ;
        RECT  0.965 3.440 2.895 3.940 ;
        RECT  0.705 2.585 0.965 3.940 ;
        RECT  0.000 3.440 0.705 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.080 1.785 3.210 2.045 ;
        RECT  2.920 1.785 3.080 2.920 ;
        RECT  2.135 2.760 2.920 2.920 ;
        RECT  2.475 0.535 2.615 0.695 ;
        RECT  2.475 2.305 2.575 2.565 ;
        RECT  2.315 0.535 2.475 2.565 ;
        RECT  1.975 0.555 2.135 2.920 ;
        RECT  1.780 0.555 1.975 0.815 ;
        RECT  1.740 2.320 1.975 2.580 ;
        RECT  1.630 1.125 1.790 2.140 ;
        RECT  1.525 1.125 1.630 1.285 ;
        RECT  1.485 1.980 1.630 2.140 ;
        RECT  1.485 2.825 1.545 3.085 ;
        RECT  1.265 1.025 1.525 1.285 ;
        RECT  1.325 1.980 1.485 3.085 ;
        RECT  1.285 1.535 1.445 1.795 ;
        RECT  1.285 2.825 1.325 3.085 ;
        RECT  0.385 1.535 1.285 1.695 ;
        RECT  0.225 0.875 0.385 2.520 ;
        RECT  0.125 0.875 0.225 1.135 ;
        RECT  0.125 2.260 0.225 2.520 ;
    END
END MX2XL

MACRO AO22X4
    CLASS CORE ;
    FOREIGN AO22X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.700 3.555 2.585 ;
        RECT  3.240 1.700 3.500 2.895 ;
        RECT  3.070 1.700 3.240 1.990 ;
        RECT  2.975 1.700 3.070 1.900 ;
        RECT  2.775 0.510 2.975 1.900 ;
        RECT  2.570 0.510 2.775 0.770 ;
        END
        ANTENNADIFFAREA     0.8126 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.460 0.365 1.990 ;
        END
        ANTENNAGATEAREA     0.2795 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.520 1.065 1.990 ;
        END
        ANTENNAGATEAREA     0.2795 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 1.290 2.175 1.795 ;
        END
        ANTENNAGATEAREA     0.2795 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.290 1.715 1.845 ;
        RECT  1.285 1.585 1.505 1.845 ;
        END
        ANTENNAGATEAREA     0.2795 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.415 -0.250 4.140 0.250 ;
        RECT  3.155 -0.250 3.415 1.135 ;
        RECT  2.255 -0.250 3.155 0.250 ;
        RECT  1.995 -0.250 2.255 0.745 ;
        RECT  0.385 -0.250 1.995 0.250 ;
        RECT  0.125 -0.250 0.385 1.155 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 3.440 4.140 3.940 ;
        RECT  3.750 2.070 4.010 3.940 ;
        RECT  2.955 3.440 3.750 3.940 ;
        RECT  2.695 2.260 2.955 3.940 ;
        RECT  0.895 3.440 2.695 3.940 ;
        RECT  0.635 2.535 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.515 1.415 2.535 1.675 ;
        RECT  2.355 0.950 2.515 2.305 ;
        RECT  2.165 2.510 2.425 3.110 ;
        RECT  1.275 0.950 2.355 1.110 ;
        RECT  1.915 2.145 2.355 2.305 ;
        RECT  1.405 2.950 2.165 3.110 ;
        RECT  1.655 2.145 1.915 2.745 ;
        RECT  1.145 2.170 1.405 3.110 ;
        RECT  1.015 0.600 1.275 1.200 ;
        RECT  0.385 2.170 1.145 2.330 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END AO22X4

MACRO AO22X2
    CLASS CORE ;
    FOREIGN AO22X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.070 0.610 3.095 2.810 ;
        RECT  2.910 0.610 3.070 2.895 ;
        RECT  2.885 0.510 2.910 2.895 ;
        RECT  2.545 0.510 2.885 0.770 ;
        RECT  2.625 2.685 2.885 2.945 ;
        END
        ANTENNADIFFAREA     0.6144 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.460 0.365 1.990 ;
        END
        ANTENNAGATEAREA     0.1339 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.525 0.985 1.885 ;
        RECT  0.635 1.525 0.795 1.990 ;
        RECT  0.585 1.700 0.635 1.990 ;
        END
        ANTENNAGATEAREA     0.1339 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.175 1.670 ;
        RECT  1.635 1.410 1.965 1.670 ;
        END
        ANTENNAGATEAREA     0.1339 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 0.440 1.500 0.760 ;
        END
        ANTENNAGATEAREA     0.1339 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 -0.250 3.220 0.250 ;
        RECT  1.945 -0.250 2.205 0.745 ;
        RECT  0.385 -0.250 1.945 0.250 ;
        RECT  0.125 -0.250 0.385 1.210 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 3.440 3.220 3.940 ;
        RECT  1.805 3.285 2.745 3.940 ;
        RECT  0.925 3.440 1.805 3.940 ;
        RECT  0.665 2.865 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.525 1.405 2.625 1.665 ;
        RECT  2.365 0.950 2.525 1.665 ;
        RECT  2.385 2.065 2.485 2.325 ;
        RECT  2.225 2.065 2.385 2.725 ;
        RECT  1.365 0.950 2.365 1.110 ;
        RECT  1.465 2.565 2.225 2.725 ;
        RECT  1.875 2.070 1.975 2.330 ;
        RECT  1.715 1.850 1.875 2.330 ;
        RECT  1.365 1.850 1.715 2.010 ;
        RECT  1.305 2.190 1.465 2.725 ;
        RECT  1.205 0.950 1.365 2.010 ;
        RECT  1.205 2.190 1.305 2.505 ;
        RECT  0.985 0.950 1.205 1.210 ;
        RECT  0.385 2.345 1.205 2.505 ;
        RECT  0.175 2.170 0.385 2.505 ;
        RECT  0.125 2.170 0.175 2.430 ;
    END
END AO22X2

MACRO AO22X1
    CLASS CORE ;
    FOREIGN AO22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 1.005 2.635 2.895 ;
        RECT  2.425 1.005 2.475 1.355 ;
        RECT  2.425 2.520 2.475 2.895 ;
        RECT  2.375 1.005 2.425 1.165 ;
        RECT  1.730 2.735 2.425 2.895 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.460 0.365 1.990 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.425 0.875 1.755 ;
        RECT  0.585 1.290 0.795 1.755 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.340 2.185 1.650 ;
        RECT  1.965 1.290 2.175 1.650 ;
        RECT  1.775 1.340 1.965 1.650 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 0.440 1.255 0.815 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.070 -0.250 2.760 0.250 ;
        RECT  1.810 -0.250 2.070 0.405 ;
        RECT  0.385 -0.250 1.810 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 3.440 2.760 3.940 ;
        RECT  1.730 3.285 2.330 3.940 ;
        RECT  0.895 3.440 1.730 3.940 ;
        RECT  0.635 2.875 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.255 0.480 2.415 0.770 ;
        RECT  2.245 1.965 2.270 2.225 ;
        RECT  1.595 0.610 2.255 0.770 ;
        RECT  2.085 1.965 2.245 2.515 ;
        RECT  1.250 2.355 2.085 2.515 ;
        RECT  1.595 2.005 1.810 2.165 ;
        RECT  1.435 0.610 1.595 2.165 ;
        RECT  0.975 0.995 1.435 1.265 ;
        RECT  1.090 1.975 1.250 2.515 ;
        RECT  0.385 2.355 1.090 2.515 ;
        RECT  0.225 2.355 0.385 2.815 ;
        RECT  0.125 2.555 0.225 2.815 ;
    END
END AO22X1

MACRO AO22XL
    CLASS CORE ;
    FOREIGN AO22XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 2.520 2.635 2.810 ;
        RECT  2.450 0.925 2.610 2.895 ;
        RECT  2.425 0.925 2.450 1.355 ;
        RECT  2.425 2.520 2.450 2.895 ;
        RECT  1.920 2.735 2.425 2.895 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.460 0.365 1.990 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.425 0.875 1.755 ;
        RECT  0.585 1.290 0.795 1.755 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.945 1.055 2.180 1.580 ;
        RECT  1.610 1.325 1.945 1.485 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.925 0.460 1.375 0.785 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.065 -0.250 2.760 0.250 ;
        RECT  1.805 -0.250 2.065 0.405 ;
        RECT  0.385 -0.250 1.805 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.180 3.440 2.760 3.940 ;
        RECT  1.920 3.285 2.180 3.940 ;
        RECT  0.895 3.440 1.920 3.940 ;
        RECT  0.635 2.875 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.245 0.470 2.405 0.745 ;
        RECT  2.245 1.955 2.270 2.215 ;
        RECT  1.750 0.585 2.245 0.745 ;
        RECT  2.085 1.955 2.245 2.555 ;
        RECT  1.300 2.395 2.085 2.555 ;
        RECT  1.600 1.665 1.760 2.215 ;
        RECT  1.590 0.585 1.750 1.145 ;
        RECT  1.215 1.665 1.600 1.825 ;
        RECT  1.215 0.985 1.590 1.145 ;
        RECT  1.040 2.005 1.300 2.555 ;
        RECT  1.055 0.985 1.215 1.825 ;
        RECT  0.975 0.985 1.055 1.255 ;
        RECT  0.385 2.395 1.040 2.555 ;
        RECT  0.125 2.395 0.385 2.795 ;
    END
END AO22XL

MACRO AO21X4
    CLASS CORE ;
    FOREIGN AO21X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.025 3.095 2.180 ;
        RECT  2.830 1.025 2.885 1.225 ;
        RECT  2.830 1.980 2.885 2.180 ;
        RECT  2.570 0.605 2.830 1.225 ;
        RECT  2.570 1.980 2.830 2.950 ;
        END
        ANTENNADIFFAREA     0.7832 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.480 1.570 1.715 1.990 ;
        RECT  1.320 1.570 1.480 1.845 ;
        END
        ANTENNAGATEAREA     0.2522 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.285 0.355 1.850 ;
        END
        ANTENNAGATEAREA     0.2795 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.580 1.035 1.840 ;
        RECT  0.775 1.290 0.795 1.840 ;
        RECT  0.610 1.290 0.775 1.740 ;
        RECT  0.585 1.290 0.610 1.580 ;
        END
        ANTENNAGATEAREA     0.2795 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.370 -0.250 3.680 0.250 ;
        RECT  3.110 -0.250 3.370 0.840 ;
        RECT  2.265 -0.250 3.110 0.250 ;
        RECT  2.005 -0.250 2.265 0.870 ;
        RECT  0.385 -0.250 2.005 0.250 ;
        RECT  1.665 0.610 2.005 0.870 ;
        RECT  0.125 -0.250 0.385 1.075 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.340 3.440 3.680 3.940 ;
        RECT  3.080 2.415 3.340 3.940 ;
        RECT  2.320 3.440 3.080 3.940 ;
        RECT  2.060 2.955 2.320 3.940 ;
        RECT  0.895 3.440 2.060 3.940 ;
        RECT  0.635 2.605 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.385 1.405 2.660 1.665 ;
        RECT  2.225 1.125 2.385 2.525 ;
        RECT  1.235 1.125 2.225 1.285 ;
        RECT  1.920 2.365 2.225 2.525 ;
        RECT  1.660 2.365 1.920 2.625 ;
        RECT  1.145 2.170 1.405 3.110 ;
        RECT  0.975 0.685 1.235 1.285 ;
        RECT  0.385 2.170 1.145 2.330 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END AO21X4

MACRO AO21X2
    CLASS CORE ;
    FOREIGN AO21X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.500 0.695 2.635 2.585 ;
        RECT  2.495 0.695 2.500 2.840 ;
        RECT  2.340 0.475 2.495 2.840 ;
        RECT  2.335 0.475 2.340 1.925 ;
        RECT  2.320 2.680 2.340 2.840 ;
        RECT  2.235 0.475 2.335 1.075 ;
        RECT  2.060 2.680 2.320 2.940 ;
        END
        ANTENNADIFFAREA     0.6130 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.665 1.700 1.715 1.990 ;
        RECT  1.505 1.475 1.665 1.990 ;
        RECT  1.290 1.475 1.505 1.735 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.390 1.415 0.465 1.675 ;
        RECT  0.125 1.100 0.390 1.675 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 0.505 1.155 0.765 ;
        RECT  0.770 0.505 0.795 1.170 ;
        RECT  0.635 0.605 0.770 1.170 ;
        RECT  0.585 0.695 0.635 1.170 ;
        END
        ANTENNAGATEAREA     0.1313 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 -0.250 2.760 0.250 ;
        RECT  1.695 -0.250 1.955 0.735 ;
        RECT  0.405 -0.250 1.695 0.250 ;
        RECT  0.145 -0.250 0.405 0.850 ;
        RECT  0.000 -0.250 0.145 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.320 3.440 2.760 3.940 ;
        RECT  1.380 3.285 2.320 3.940 ;
        RECT  0.895 3.440 1.380 3.940 ;
        RECT  0.635 2.260 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.895 1.115 2.055 2.430 ;
        RECT  1.380 1.115 1.895 1.275 ;
        RECT  1.655 2.170 1.895 2.430 ;
        RECT  1.305 2.165 1.405 2.425 ;
        RECT  1.120 1.015 1.380 1.275 ;
        RECT  1.145 1.920 1.305 2.425 ;
        RECT  0.385 1.920 1.145 2.080 ;
        RECT  0.125 1.920 0.385 2.555 ;
    END
END AO21X2

MACRO AO21X1
    CLASS CORE ;
    FOREIGN AO21X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.135 1.515 2.175 1.990 ;
        RECT  2.125 1.515 2.135 2.810 ;
        RECT  1.975 1.035 2.125 2.810 ;
        RECT  1.965 1.035 1.975 1.990 ;
        RECT  1.875 2.650 1.975 2.810 ;
        RECT  1.615 2.650 1.875 2.910 ;
        END
        ANTENNADIFFAREA     0.3398 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.565 1.425 1.990 ;
        END
        ANTENNAGATEAREA     0.0624 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.240 0.445 1.665 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 2.520 1.165 2.810 ;
        END
        ANTENNAGATEAREA     0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 -0.250 2.300 0.250 ;
        RECT  1.295 -0.250 1.555 0.405 ;
        RECT  0.385 -0.250 1.295 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.870 3.440 2.300 3.940 ;
        RECT  0.930 3.285 1.870 3.940 ;
        RECT  0.000 3.440 0.930 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.765 0.545 1.995 0.805 ;
        RECT  1.765 2.140 1.795 2.400 ;
        RECT  1.735 0.545 1.765 2.400 ;
        RECT  1.605 0.645 1.735 2.400 ;
        RECT  1.125 1.135 1.605 1.295 ;
        RECT  0.385 2.170 1.335 2.330 ;
        RECT  0.865 1.035 1.125 1.295 ;
        RECT  0.125 2.120 0.385 2.380 ;
    END
END AO21X1

MACRO AO21XL
    CLASS CORE ;
    FOREIGN AO21XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.135 1.515 2.175 1.990 ;
        RECT  2.125 1.515 2.135 2.810 ;
        RECT  1.975 1.030 2.125 2.810 ;
        RECT  1.965 1.030 1.975 1.990 ;
        RECT  1.875 2.650 1.975 2.810 ;
        RECT  1.615 2.650 1.875 2.910 ;
        END
        ANTENNADIFFAREA     0.2188 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.565 1.425 1.990 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.240 0.445 1.665 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 2.520 1.165 2.810 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 -0.250 2.300 0.250 ;
        RECT  1.295 -0.250 1.555 0.405 ;
        RECT  0.385 -0.250 1.295 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.875 3.440 2.300 3.940 ;
        RECT  0.935 3.285 1.875 3.940 ;
        RECT  0.000 3.440 0.935 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.785 0.545 1.995 0.805 ;
        RECT  1.785 2.120 1.795 2.380 ;
        RECT  1.735 0.545 1.785 2.380 ;
        RECT  1.625 0.645 1.735 2.380 ;
        RECT  1.615 0.645 1.625 1.295 ;
        RECT  1.125 1.135 1.615 1.295 ;
        RECT  0.385 2.170 1.335 2.330 ;
        RECT  0.865 1.035 1.125 1.295 ;
        RECT  0.125 2.120 0.385 2.380 ;
    END
END AO21XL

MACRO AOI2BB2X4
    CLASS CORE ;
    FOREIGN AOI2BB2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.515 0.615 6.775 0.875 ;
        RECT  4.280 0.635 6.515 0.875 ;
        RECT  4.040 0.635 4.280 1.285 ;
        RECT  2.875 1.045 4.040 1.285 ;
        RECT  3.085 2.015 3.345 2.725 ;
        RECT  2.650 2.015 3.085 2.255 ;
        RECT  2.650 0.495 2.875 1.285 ;
        RECT  2.615 0.495 2.650 2.255 ;
        RECT  2.410 1.045 2.615 2.255 ;
        RECT  2.325 2.015 2.410 2.255 ;
        RECT  2.065 2.015 2.325 3.035 ;
        RECT  1.965 2.335 2.065 2.585 ;
        END
        ANTENNADIFFAREA     1.6408 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.735 1.745 5.995 2.005 ;
        RECT  5.380 1.845 5.735 2.005 ;
        RECT  5.120 1.395 5.380 2.005 ;
        RECT  4.015 1.845 5.120 2.005 ;
        RECT  3.995 1.700 4.015 2.005 ;
        RECT  3.805 1.560 3.995 2.005 ;
        RECT  3.735 1.560 3.805 1.820 ;
        END
        ANTENNAGATEAREA     0.6630 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.505 1.265 6.605 1.525 ;
        RECT  6.345 1.055 6.505 1.525 ;
        RECT  4.935 1.055 6.345 1.215 ;
        RECT  4.775 1.055 4.935 1.665 ;
        RECT  4.725 1.290 4.775 1.665 ;
        RECT  4.460 1.405 4.725 1.665 ;
        END
        ANTENNAGATEAREA     0.7098 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.575 1.750 1.835 ;
        RECT  1.650 1.575 1.715 2.810 ;
        RECT  1.490 1.575 1.650 3.025 ;
        RECT  0.370 2.865 1.490 3.025 ;
        RECT  0.210 1.575 0.370 3.025 ;
        RECT  0.125 1.575 0.210 2.585 ;
        RECT  0.110 1.575 0.125 1.835 ;
        END
        ANTENNAGATEAREA     0.3003 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.455 0.930 1.990 ;
        END
        ANTENNAGATEAREA     0.3003 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.920 -0.250 6.900 0.250 ;
        RECT  5.320 -0.250 5.920 0.405 ;
        RECT  3.815 -0.250 5.320 0.250 ;
        RECT  3.215 -0.250 3.815 0.825 ;
        RECT  2.335 -0.250 3.215 0.250 ;
        RECT  1.735 -0.250 2.335 0.825 ;
        RECT  0.910 -0.250 1.735 0.250 ;
        RECT  0.650 -0.250 0.910 1.165 ;
        RECT  0.000 -0.250 0.650 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.375 3.440 6.900 3.940 ;
        RECT  6.115 3.285 6.375 3.940 ;
        RECT  5.315 3.440 6.115 3.940 ;
        RECT  5.055 2.645 5.315 3.940 ;
        RECT  4.255 3.440 5.055 3.940 ;
        RECT  3.995 3.285 4.255 3.940 ;
        RECT  1.810 3.440 3.995 3.940 ;
        RECT  1.550 3.285 1.810 3.940 ;
        RECT  0.385 3.440 1.550 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.515 1.975 6.775 2.915 ;
        RECT  5.825 2.255 6.515 2.415 ;
        RECT  5.565 2.255 5.825 2.915 ;
        RECT  4.805 2.255 5.565 2.415 ;
        RECT  4.545 2.255 4.805 3.195 ;
        RECT  3.855 2.255 4.545 2.415 ;
        RECT  3.755 2.255 3.855 2.915 ;
        RECT  3.595 2.255 3.755 3.085 ;
        RECT  2.835 2.925 3.595 3.085 ;
        RECT  2.675 2.435 2.835 3.085 ;
        RECT  2.575 2.435 2.675 3.035 ;
        RECT  2.130 1.575 2.230 1.835 ;
        RECT  1.970 1.235 2.130 1.835 ;
        RECT  1.450 1.235 1.970 1.395 ;
        RECT  1.270 0.595 1.450 1.395 ;
        RECT  1.190 0.595 1.270 2.470 ;
        RECT  1.110 1.230 1.190 2.470 ;
        RECT  0.840 2.210 1.110 2.470 ;
    END
END AOI2BB2X4

MACRO AOI2BB2X2
    CLASS CORE ;
    FOREIGN AOI2BB2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.985 2.110 4.015 2.400 ;
        RECT  3.825 0.925 3.985 2.400 ;
        RECT  2.120 0.925 3.825 1.085 ;
        RECT  3.805 2.110 3.825 2.400 ;
        RECT  3.045 2.170 3.805 2.330 ;
        RECT  2.785 2.020 3.045 2.620 ;
        END
        ANTENNADIFFAREA     0.7789 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.265 3.645 1.925 ;
        RECT  3.345 1.265 3.555 1.990 ;
        RECT  2.265 1.265 3.345 1.425 ;
        RECT  2.105 1.265 2.265 2.145 ;
        RECT  1.300 1.985 2.105 2.145 ;
        RECT  1.090 1.760 1.300 2.145 ;
        END
        ANTENNAGATEAREA     0.3536 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.770 0.470 4.030 0.745 ;
        RECT  1.925 0.585 3.770 0.745 ;
        RECT  1.765 0.585 1.925 1.800 ;
        RECT  1.505 1.290 1.765 1.800 ;
        END
        ANTENNAGATEAREA     0.3536 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.865 1.270 1.325 1.580 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.270 0.345 1.990 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.920 -0.250 4.140 0.250 ;
        RECT  2.660 -0.250 2.920 0.405 ;
        RECT  1.500 -0.250 2.660 0.250 ;
        RECT  1.240 -0.250 1.500 1.085 ;
        RECT  0.385 -0.250 1.240 0.250 ;
        RECT  0.335 -0.250 0.385 0.405 ;
        RECT  0.175 -0.250 0.335 1.080 ;
        RECT  0.125 -0.250 0.175 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 3.285 4.015 3.940 ;
        RECT  2.055 3.440 3.755 3.940 ;
        RECT  1.795 3.285 2.055 3.940 ;
        RECT  1.250 3.440 1.795 3.940 ;
        RECT  0.990 3.285 1.250 3.940 ;
        RECT  0.000 3.440 0.990 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.485 2.520 3.585 2.780 ;
        RECT  3.325 2.520 3.485 2.960 ;
        RECT  2.645 2.800 3.325 2.960 ;
        RECT  2.605 1.605 2.810 1.765 ;
        RECT  2.385 2.800 2.645 3.220 ;
        RECT  2.445 1.605 2.605 2.485 ;
        RECT  0.685 2.325 2.445 2.485 ;
        RECT  1.650 2.800 2.385 2.960 ;
        RECT  1.390 2.665 1.650 2.960 ;
        RECT  0.685 0.830 0.905 1.090 ;
        RECT  0.590 0.830 0.685 2.485 ;
        RECT  0.525 0.830 0.590 2.575 ;
        RECT  0.385 2.250 0.525 2.575 ;
        RECT  0.125 2.250 0.385 2.850 ;
    END
END AOI2BB2X2

MACRO AOI2BB2X1
    CLASS CORE ;
    FOREIGN AOI2BB2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.105 2.635 2.855 ;
        RECT  2.425 1.005 2.585 2.855 ;
        RECT  2.110 1.005 2.425 1.165 ;
        RECT  2.375 2.255 2.425 2.855 ;
        RECT  1.850 0.875 2.110 1.165 ;
        END
        ANTENNADIFFAREA     0.4376 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 2.930 1.255 3.220 ;
        RECT  0.725 2.945 1.045 3.105 ;
        RECT  0.465 2.845 0.725 3.105 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 2.110 2.175 2.400 ;
        RECT  1.815 2.110 1.965 2.270 ;
        RECT  1.650 1.830 1.815 2.270 ;
        RECT  1.555 1.830 1.650 2.090 ;
        END
        ANTENNAGATEAREA     0.1651 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.175 1.430 0.335 2.400 ;
        RECT  0.125 1.925 0.175 2.400 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.925 1.775 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 -0.250 2.760 0.250 ;
        RECT  2.375 -0.250 2.635 0.405 ;
        RECT  1.385 -0.250 2.375 0.250 ;
        RECT  1.125 -0.250 1.385 0.405 ;
        RECT  0.385 -0.250 1.125 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.705 3.440 2.760 3.940 ;
        RECT  1.445 3.285 1.705 3.940 ;
        RECT  0.385 3.440 1.445 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.085 1.345 2.245 1.625 ;
        RECT  1.865 2.580 2.125 2.910 ;
        RECT  1.265 1.345 2.085 1.505 ;
        RECT  0.905 2.580 1.865 2.740 ;
        RECT  1.105 0.950 1.265 2.155 ;
        RECT  0.820 0.950 1.105 1.110 ;
        RECT  1.095 1.970 1.105 2.155 ;
        RECT  0.835 1.970 1.095 2.230 ;
        RECT  0.560 0.850 0.820 1.110 ;
    END
END AOI2BB2X1

MACRO AOI2BB2XL
    CLASS CORE ;
    FOREIGN AOI2BB2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.615 1.515 2.635 2.810 ;
        RECT  2.515 1.515 2.615 2.945 ;
        RECT  2.355 1.095 2.515 2.945 ;
        RECT  2.060 1.095 2.355 1.255 ;
        RECT  1.900 0.985 2.060 1.255 ;
        END
        ANTENNADIFFAREA     0.2738 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.605 1.290 1.715 1.580 ;
        RECT  1.505 1.290 1.605 1.945 ;
        RECT  1.445 1.355 1.505 1.945 ;
        END
        ANTENNAGATEAREA     0.0975 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.990 1.700 2.175 2.325 ;
        RECT  1.965 1.700 1.990 2.425 ;
        RECT  1.680 2.165 1.965 2.425 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.365 0.405 1.625 ;
        RECT  0.145 1.365 0.335 2.400 ;
        RECT  0.125 1.515 0.145 2.400 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.880 1.775 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.540 -0.250 2.760 0.250 ;
        RECT  2.280 -0.250 2.540 0.405 ;
        RECT  1.400 -0.250 2.280 0.250 ;
        RECT  1.140 -0.250 1.400 0.405 ;
        RECT  0.390 -0.250 1.140 0.250 ;
        RECT  0.130 -0.250 0.390 0.405 ;
        RECT  0.000 -0.250 0.130 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 3.440 2.760 3.940 ;
        RECT  1.245 2.945 1.505 3.940 ;
        RECT  0.390 3.440 1.245 3.940 ;
        RECT  0.130 2.605 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.990 0.585 2.250 0.775 ;
        RECT  1.845 2.605 2.105 2.945 ;
        RECT  1.265 0.585 1.990 0.745 ;
        RECT  0.900 2.605 1.845 2.765 ;
        RECT  1.105 0.585 1.265 2.115 ;
        RECT  0.820 0.585 1.105 0.745 ;
        RECT  1.100 1.955 1.105 2.115 ;
        RECT  0.840 1.955 1.100 2.215 ;
        RECT  0.640 2.605 0.900 2.885 ;
        RECT  0.660 0.585 0.820 1.110 ;
        RECT  0.560 0.950 0.660 1.110 ;
    END
END AOI2BB2XL

MACRO AOI2BB1X4
    CLASS CORE ;
    FOREIGN AOI2BB1X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 1.515 4.475 3.215 ;
        RECT  4.215 0.935 4.385 3.215 ;
        RECT  4.145 0.935 4.215 2.435 ;
        RECT  4.015 0.935 4.145 1.175 ;
        RECT  3.990 2.110 4.145 2.435 ;
        RECT  3.965 0.695 4.015 1.175 ;
        RECT  2.835 2.195 3.990 2.435 ;
        RECT  3.705 0.575 3.965 1.175 ;
        RECT  2.940 0.935 3.705 1.175 ;
        RECT  2.680 0.495 2.940 1.175 ;
        RECT  2.575 2.195 2.835 3.190 ;
        RECT  2.425 2.745 2.575 3.190 ;
        END
        ANTENNADIFFAREA     1.4506 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.225 1.750 3.485 2.010 ;
        RECT  3.095 1.750 3.225 1.990 ;
        RECT  2.885 1.700 3.095 1.990 ;
        END
        ANTENNAGATEAREA     0.6552 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.585 1.790 1.845 ;
        RECT  1.665 1.585 1.715 2.400 ;
        RECT  1.505 1.585 1.665 2.675 ;
        RECT  1.435 2.515 1.505 2.675 ;
        RECT  1.275 2.515 1.435 2.770 ;
        RECT  0.370 2.610 1.275 2.770 ;
        RECT  0.125 1.575 0.370 2.770 ;
        RECT  0.110 1.575 0.125 1.835 ;
        END
        ANTENNAGATEAREA     0.3003 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.665 1.575 0.925 1.990 ;
        RECT  0.585 1.700 0.665 1.990 ;
        END
        ANTENNAGATEAREA     0.3003 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 -0.250 4.600 0.250 ;
        RECT  4.215 -0.250 4.475 0.755 ;
        RECT  3.455 -0.250 4.215 0.250 ;
        RECT  3.195 -0.250 3.455 0.755 ;
        RECT  2.430 -0.250 3.195 0.250 ;
        RECT  2.170 -0.250 2.430 1.045 ;
        RECT  1.110 -0.250 2.170 0.250 ;
        RECT  0.850 -0.250 1.110 1.000 ;
        RECT  0.000 -0.250 0.850 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.655 3.440 4.600 3.940 ;
        RECT  3.395 2.615 3.655 3.940 ;
        RECT  1.975 3.440 3.395 3.940 ;
        RECT  1.715 2.895 1.975 3.940 ;
        RECT  0.385 3.440 1.715 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.705 1.355 3.965 1.705 ;
        RECT  2.665 1.355 3.705 1.515 ;
        RECT  2.405 1.355 2.665 1.995 ;
        RECT  2.215 1.355 2.405 1.515 ;
        RECT  2.055 1.245 2.215 1.515 ;
        RECT  1.620 1.245 2.055 1.405 ;
        RECT  1.360 0.695 1.620 1.405 ;
        RECT  1.325 1.235 1.360 1.405 ;
        RECT  1.165 1.235 1.325 2.330 ;
        RECT  0.600 1.235 1.165 1.395 ;
        RECT  1.095 2.170 1.165 2.330 ;
        RECT  0.835 2.170 1.095 2.430 ;
        RECT  0.340 0.695 0.600 1.395 ;
    END
END AOI2BB1X4

MACRO AOI2BB1X2
    CLASS CORE ;
    FOREIGN AOI2BB1X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.890 1.035 1.925 2.270 ;
        RECT  1.765 1.035 1.890 2.715 ;
        RECT  1.630 2.110 1.765 2.715 ;
        RECT  1.505 2.110 1.630 2.400 ;
        END
        ANTENNADIFFAREA     0.6384 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.440 1.700 2.635 1.990 ;
        RECT  2.425 0.690 2.440 1.990 ;
        RECT  2.280 0.690 2.425 1.985 ;
        RECT  1.555 0.690 2.280 0.850 ;
        RECT  1.395 0.690 1.555 1.665 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.715 1.585 0.875 2.400 ;
        RECT  0.585 2.110 0.715 2.400 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.490 0.445 1.750 ;
        RECT  0.125 1.490 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.515 -0.250 2.760 0.250 ;
        RECT  2.255 -0.250 2.515 0.405 ;
        RECT  1.435 -0.250 2.255 0.250 ;
        RECT  1.175 -0.250 1.435 0.405 ;
        RECT  0.385 -0.250 1.175 0.250 ;
        RECT  0.125 -0.250 0.385 1.065 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.600 3.440 2.760 3.940 ;
        RECT  2.340 3.285 2.600 3.940 ;
        RECT  0.985 3.440 2.340 3.940 ;
        RECT  0.725 3.285 0.985 3.940 ;
        RECT  0.000 3.440 0.725 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.800 2.945 2.060 3.215 ;
        RECT  1.215 2.945 1.800 3.105 ;
        RECT  1.055 0.955 1.215 3.105 ;
        RECT  0.895 0.955 1.055 1.115 ;
        RECT  0.385 2.945 1.055 3.105 ;
        RECT  0.635 0.855 0.895 1.115 ;
        RECT  0.125 2.945 0.385 3.255 ;
    END
END AOI2BB1X2

MACRO AOI2BB1X1
    CLASS CORE ;
    FOREIGN AOI2BB1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.075 2.200 2.175 ;
        RECT  2.125 1.075 2.175 2.585 ;
        RECT  2.040 1.075 2.125 2.930 ;
        RECT  1.770 1.075 2.040 1.235 ;
        RECT  2.015 2.000 2.040 2.930 ;
        RECT  1.965 2.110 2.015 2.930 ;
        RECT  1.865 2.230 1.965 2.930 ;
        RECT  1.510 0.975 1.770 1.235 ;
        END
        ANTENNADIFFAREA     0.4830 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.760 1.345 2.400 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.640 0.795 2.400 ;
        RECT  0.535 1.640 0.585 1.900 ;
        END
        ANTENNAGATEAREA     0.0741 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.120 0.370 2.380 ;
        RECT  0.125 1.700 0.335 2.380 ;
        RECT  0.110 2.120 0.125 2.380 ;
        END
        ANTENNAGATEAREA     0.0741 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.170 -0.250 2.300 0.250 ;
        RECT  1.230 -0.250 2.170 0.405 ;
        RECT  0.920 -0.250 1.230 0.250 ;
        RECT  0.660 -0.250 0.920 0.405 ;
        RECT  0.000 -0.250 0.660 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.095 3.440 2.300 3.940 ;
        RECT  0.835 3.285 1.095 3.940 ;
        RECT  0.000 3.440 0.835 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.685 1.415 1.860 1.675 ;
        RECT  1.525 1.415 1.685 2.920 ;
        RECT  1.135 1.415 1.525 1.575 ;
        RECT  0.385 2.760 1.525 2.920 ;
        RECT  0.975 1.135 1.135 1.575 ;
        RECT  0.580 1.135 0.975 1.295 ;
        RECT  0.320 1.035 0.580 1.295 ;
        RECT  0.125 2.580 0.385 2.920 ;
    END
END AOI2BB1X1

MACRO AOI2BB1XL
    CLASS CORE ;
    FOREIGN AOI2BB1XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.015 1.135 2.175 2.525 ;
        RECT  1.980 1.135 2.015 1.295 ;
        RECT  1.965 2.110 2.015 2.525 ;
        RECT  1.720 1.035 1.980 1.295 ;
        RECT  1.865 2.265 1.965 2.525 ;
        END
        ANTENNADIFFAREA     0.3330 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.815 1.345 2.075 ;
        RECT  1.085 1.815 1.255 2.400 ;
        RECT  1.045 2.110 1.085 2.400 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.495 0.865 1.755 ;
        RECT  0.605 1.495 0.795 2.400 ;
        RECT  0.585 1.755 0.605 2.400 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.490 0.370 2.005 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.170 -0.250 2.300 0.250 ;
        RECT  1.230 -0.250 2.170 0.405 ;
        RECT  0.920 -0.250 1.230 0.250 ;
        RECT  0.660 -0.250 0.920 0.405 ;
        RECT  0.000 -0.250 0.660 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 3.440 2.300 3.940 ;
        RECT  0.975 2.945 1.235 3.940 ;
        RECT  0.000 3.440 0.975 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.685 1.475 1.820 1.735 ;
        RECT  1.525 1.475 1.685 2.740 ;
        RECT  1.320 1.475 1.525 1.635 ;
        RECT  0.385 2.580 1.525 2.740 ;
        RECT  1.160 1.135 1.320 1.635 ;
        RECT  0.580 1.135 1.160 1.295 ;
        RECT  0.320 1.035 0.580 1.295 ;
        RECT  0.225 2.185 0.385 2.740 ;
        RECT  0.125 2.185 0.225 2.445 ;
    END
END AOI2BB1XL

MACRO AOI33X4
    CLASS CORE ;
    FOREIGN AOI33X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.915 1.290 4.935 2.175 ;
        RECT  4.715 0.975 4.915 2.325 ;
        RECT  4.475 0.975 4.715 1.175 ;
        RECT  4.475 2.125 4.715 2.325 ;
        RECT  4.425 0.695 4.475 1.175 ;
        RECT  4.420 2.125 4.475 2.585 ;
        RECT  4.165 0.575 4.425 1.175 ;
        RECT  4.160 2.125 4.420 3.065 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.215 0.370 1.990 ;
        RECT  0.110 1.215 0.125 1.475 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.525 0.925 1.785 ;
        RECT  0.635 0.880 0.795 1.785 ;
        RECT  0.585 0.880 0.635 1.355 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 1.025 1.375 1.285 ;
        RECT  1.105 1.025 1.265 2.400 ;
        RECT  1.045 2.110 1.105 2.400 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.700 3.095 1.990 ;
        RECT  2.765 1.700 2.885 1.860 ;
        RECT  2.605 1.285 2.765 1.860 ;
        RECT  2.505 1.285 2.605 1.545 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.080 2.635 2.400 ;
        RECT  2.285 2.080 2.425 2.240 ;
        RECT  2.125 1.765 2.285 2.240 ;
        RECT  2.025 1.765 2.125 2.025 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.805 1.290 2.175 1.580 ;
        RECT  1.645 1.290 1.805 2.095 ;
        RECT  1.545 1.835 1.645 2.095 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 -0.250 5.060 0.250 ;
        RECT  4.675 -0.250 4.935 0.755 ;
        RECT  3.860 -0.250 4.675 0.250 ;
        RECT  3.700 -0.250 3.860 0.815 ;
        RECT  2.680 -0.250 3.700 0.250 ;
        RECT  2.420 -0.250 2.680 0.765 ;
        RECT  0.385 -0.250 2.420 0.250 ;
        RECT  0.125 -0.250 0.385 0.795 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 3.440 5.060 3.940 ;
        RECT  4.675 2.595 4.935 3.940 ;
        RECT  3.870 3.440 4.675 3.940 ;
        RECT  3.610 3.285 3.870 3.940 ;
        RECT  1.115 3.440 3.610 3.940 ;
        RECT  0.855 3.285 1.115 3.940 ;
        RECT  0.385 3.440 0.855 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.780 1.415 4.435 1.675 ;
        RECT  3.620 0.995 3.780 3.090 ;
        RECT  3.520 0.995 3.620 1.155 ;
        RECT  3.360 2.930 3.620 3.090 ;
        RECT  3.360 0.605 3.520 1.155 ;
        RECT  3.275 1.335 3.435 2.390 ;
        RECT  3.140 0.605 3.360 0.765 ;
        RECT  3.100 2.930 3.360 3.190 ;
        RECT  3.165 1.335 3.275 1.495 ;
        RECT  3.010 2.230 3.275 2.390 ;
        RECT  3.005 0.945 3.165 1.495 ;
        RECT  2.850 2.230 3.010 2.740 ;
        RECT  2.240 0.945 3.005 1.105 ;
        RECT  2.110 2.580 2.850 2.740 ;
        RECT  2.400 2.945 2.660 3.210 ;
        RECT  1.625 2.945 2.400 3.105 ;
        RECT  2.080 0.655 2.240 1.105 ;
        RECT  1.850 2.420 2.110 2.740 ;
        RECT  1.545 0.655 2.080 0.815 ;
        RECT  1.365 2.945 1.625 3.210 ;
        RECT  1.285 0.555 1.545 0.815 ;
        RECT  0.755 2.945 1.365 3.105 ;
        RECT  0.495 2.725 0.755 3.105 ;
    END
END AOI33X4

MACRO AOI33X2
    CLASS CORE ;
    FOREIGN AOI33X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.785 0.595 5.855 2.585 ;
        RECT  5.695 0.595 5.785 2.835 ;
        RECT  4.365 0.595 5.695 0.755 ;
        RECT  5.625 1.700 5.695 2.835 ;
        RECT  5.525 2.170 5.625 2.835 ;
        RECT  4.765 2.170 5.525 2.330 ;
        RECT  4.505 2.170 4.765 2.835 ;
        RECT  3.745 2.170 4.505 2.330 ;
        RECT  3.990 0.495 4.365 0.755 ;
        RECT  1.685 0.595 3.990 0.755 ;
        RECT  3.485 2.170 3.745 2.835 ;
        RECT  1.425 0.495 1.685 0.755 ;
        END
        ANTENNADIFFAREA     1.4592 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.795 1.795 2.935 1.955 ;
        RECT  2.635 1.795 2.795 2.330 ;
        RECT  0.340 2.170 2.635 2.330 ;
        RECT  0.340 1.235 0.555 1.495 ;
        RECT  0.180 1.235 0.340 2.330 ;
        RECT  0.125 1.515 0.180 1.990 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 1.545 2.455 1.805 ;
        RECT  2.195 0.990 2.355 1.805 ;
        RECT  1.035 0.990 2.195 1.150 ;
        RECT  2.175 1.580 2.195 1.805 ;
        RECT  1.965 1.580 2.175 1.990 ;
        RECT  0.875 0.990 1.035 1.805 ;
        RECT  0.775 1.545 0.875 1.805 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.515 1.700 1.715 1.990 ;
        RECT  1.355 1.330 1.515 1.990 ;
        RECT  1.255 1.330 1.355 1.590 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 1.225 5.495 1.485 ;
        RECT  5.235 0.950 5.395 1.485 ;
        RECT  3.390 0.950 5.235 1.110 ;
        RECT  3.230 0.950 3.390 1.540 ;
        RECT  3.095 1.280 3.230 1.540 ;
        RECT  2.885 1.290 3.095 1.580 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.915 1.545 5.015 1.805 ;
        RECT  4.755 1.545 4.915 1.990 ;
        RECT  4.015 1.830 4.755 1.990 ;
        RECT  3.805 1.700 4.015 1.990 ;
        RECT  3.625 1.730 3.805 1.990 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.195 1.290 4.575 1.650 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.525 -0.250 6.440 0.250 ;
        RECT  5.265 -0.250 5.525 0.405 ;
        RECT  3.185 -0.250 5.265 0.250 ;
        RECT  2.585 -0.250 3.185 0.405 ;
        RECT  0.525 -0.250 2.585 0.250 ;
        RECT  0.265 -0.250 0.525 0.795 ;
        RECT  0.000 -0.250 0.265 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.685 3.440 6.440 3.940 ;
        RECT  2.425 3.285 2.685 3.940 ;
        RECT  1.735 3.440 2.425 3.940 ;
        RECT  1.475 3.285 1.735 3.940 ;
        RECT  0.785 3.440 1.475 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.195 2.220 6.295 2.820 ;
        RECT  6.035 2.220 6.195 3.175 ;
        RECT  5.275 3.015 6.035 3.175 ;
        RECT  5.015 2.510 5.275 3.175 ;
        RECT  4.255 3.015 5.015 3.175 ;
        RECT  3.995 2.510 4.255 3.175 ;
        RECT  3.235 3.015 3.995 3.175 ;
        RECT  2.975 2.435 3.235 3.175 ;
        RECT  2.285 2.510 2.975 2.670 ;
        RECT  2.025 2.510 2.285 2.770 ;
        RECT  1.335 2.510 2.025 2.670 ;
        RECT  1.075 2.510 1.335 2.770 ;
        RECT  0.385 2.510 1.075 2.670 ;
        RECT  0.125 2.510 0.385 2.770 ;
    END
END AOI33X2

MACRO AOI33X1
    CLASS CORE ;
    FOREIGN AOI33X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.510 1.105 3.555 2.585 ;
        RECT  3.505 1.105 3.510 2.775 ;
        RECT  3.345 1.000 3.505 2.775 ;
        RECT  2.670 1.000 3.345 1.160 ;
        RECT  3.250 2.175 3.345 2.775 ;
        RECT  2.490 2.220 3.250 2.380 ;
        RECT  2.510 0.950 2.670 1.160 ;
        RECT  1.745 0.950 2.510 1.110 ;
        RECT  2.230 2.220 2.490 2.495 ;
        RECT  1.485 0.560 1.745 1.110 ;
        END
        ANTENNADIFFAREA     1.1676 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.340 0.405 1.600 ;
        RECT  0.145 1.340 0.335 1.990 ;
        RECT  0.125 1.700 0.145 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.630 1.040 1.890 ;
        RECT  0.635 1.290 0.795 1.890 ;
        RECT  0.585 1.290 0.635 1.765 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.620 1.640 1.880 ;
        RECT  1.380 1.290 1.540 1.880 ;
        RECT  1.255 1.290 1.380 1.450 ;
        RECT  1.095 0.880 1.255 1.450 ;
        RECT  1.045 0.880 1.095 1.170 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.100 1.340 3.150 1.600 ;
        RECT  3.095 1.340 3.100 1.925 ;
        RECT  2.890 1.340 3.095 1.990 ;
        RECT  2.885 1.700 2.890 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 1.515 2.635 2.040 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.860 1.515 2.175 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.110 -0.250 3.680 0.250 ;
        RECT  2.850 -0.250 3.110 0.820 ;
        RECT  0.390 -0.250 2.850 0.250 ;
        RECT  0.130 -0.250 0.390 1.160 ;
        RECT  0.000 -0.250 0.130 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.440 3.440 3.680 3.940 ;
        RECT  1.180 2.605 1.440 3.940 ;
        RECT  0.390 3.440 1.180 3.940 ;
        RECT  0.130 2.220 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.740 2.560 3.000 2.835 ;
        RECT  1.980 2.675 2.740 2.835 ;
        RECT  1.720 2.170 1.980 2.835 ;
        RECT  0.900 2.170 1.720 2.330 ;
        RECT  0.640 2.170 0.900 2.770 ;
    END
END AOI33X1

MACRO AOI33XL
    CLASS CORE ;
    FOREIGN AOI33XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.525 2.110 3.555 2.570 ;
        RECT  3.365 0.950 3.525 2.570 ;
        RECT  1.990 0.950 3.365 1.110 ;
        RECT  3.295 2.040 3.365 2.570 ;
        RECT  2.535 2.040 3.295 2.200 ;
        RECT  2.375 2.040 2.535 2.570 ;
        RECT  2.275 2.310 2.375 2.570 ;
        RECT  1.625 0.850 1.990 1.110 ;
        END
        ANTENNADIFFAREA     0.5640 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 1.760 0.520 2.020 ;
        RECT  0.245 1.290 0.405 2.020 ;
        RECT  0.125 1.290 0.245 1.765 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.865 1.790 1.125 2.050 ;
        RECT  0.705 1.290 0.865 2.050 ;
        RECT  0.585 1.290 0.705 1.580 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.535 1.600 1.635 1.860 ;
        RECT  1.375 1.420 1.535 1.860 ;
        RECT  1.255 1.420 1.375 1.580 ;
        RECT  1.045 1.290 1.255 1.580 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 1.540 3.185 1.860 ;
        RECT  2.885 1.290 3.095 1.860 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.540 2.655 1.860 ;
        RECT  2.425 1.290 2.635 1.860 ;
        RECT  2.395 1.540 2.425 1.860 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 1.290 2.175 1.765 ;
        RECT  1.965 1.290 2.145 1.860 ;
        RECT  1.885 1.600 1.965 1.860 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.135 -0.250 3.680 0.250 ;
        RECT  2.875 -0.250 3.135 0.745 ;
        RECT  0.615 -0.250 2.875 0.250 ;
        RECT  0.355 -0.250 0.615 0.795 ;
        RECT  0.000 -0.250 0.355 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 3.440 3.680 3.940 ;
        RECT  1.175 2.605 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.380 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.945 2.380 3.045 2.640 ;
        RECT  2.785 2.380 2.945 2.910 ;
        RECT  2.025 2.750 2.785 2.910 ;
        RECT  1.865 2.265 2.025 2.910 ;
        RECT  1.765 2.265 1.865 2.570 ;
        RECT  0.895 2.265 1.765 2.425 ;
        RECT  0.635 2.265 0.895 2.570 ;
    END
END AOI33XL

MACRO AOI32X4
    CLASS CORE ;
    FOREIGN AOI32X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 1.515 4.475 2.400 ;
        RECT  4.265 1.095 4.465 2.400 ;
        RECT  3.965 1.095 4.265 1.295 ;
        RECT  4.015 2.090 4.265 2.400 ;
        RECT  3.965 2.090 4.015 2.585 ;
        RECT  3.705 0.695 3.965 1.295 ;
        RECT  3.705 2.090 3.965 3.030 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 0.995 2.635 1.580 ;
        RECT  2.365 0.995 2.425 1.515 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 1.080 2.175 1.580 ;
        END
        ANTENNAGATEAREA     0.1079 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.295 0.445 1.555 ;
        RECT  0.150 1.295 0.335 2.400 ;
        RECT  0.125 1.515 0.150 2.400 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.585 0.925 1.845 ;
        RECT  0.665 1.585 0.795 2.400 ;
        RECT  0.635 1.635 0.665 2.400 ;
        RECT  0.585 1.925 0.635 2.400 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 1.335 1.355 1.595 ;
        RECT  1.255 1.335 1.265 2.335 ;
        RECT  1.105 1.335 1.255 2.400 ;
        RECT  1.045 2.110 1.105 2.400 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 -0.250 4.600 0.250 ;
        RECT  4.215 -0.250 4.475 0.815 ;
        RECT  3.455 -0.250 4.215 0.250 ;
        RECT  3.195 -0.250 3.455 0.815 ;
        RECT  2.370 -0.250 3.195 0.250 ;
        RECT  2.110 -0.250 2.370 0.815 ;
        RECT  0.385 -0.250 2.110 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 3.440 4.600 3.940 ;
        RECT  4.215 2.595 4.475 3.940 ;
        RECT  3.415 3.440 4.215 3.940 ;
        RECT  3.155 3.285 3.415 3.940 ;
        RECT  1.115 3.440 3.155 3.940 ;
        RECT  0.855 3.285 1.115 3.940 ;
        RECT  0.385 3.440 0.855 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.470 1.570 3.970 1.830 ;
        RECT  3.310 0.995 3.470 2.820 ;
        RECT  3.010 0.995 3.310 1.155 ;
        RECT  2.955 2.660 3.310 2.820 ;
        RECT  2.870 1.580 3.130 1.920 ;
        RECT  2.850 0.555 3.010 1.155 ;
        RECT  2.795 2.660 2.955 3.200 ;
        RECT  2.005 1.760 2.870 1.920 ;
        RECT  2.685 0.555 2.850 0.815 ;
        RECT  2.695 2.940 2.795 3.200 ;
        RECT  2.515 2.240 2.615 2.500 ;
        RECT  2.355 2.240 2.515 2.985 ;
        RECT  1.625 2.825 2.355 2.985 ;
        RECT  2.005 2.335 2.105 2.595 ;
        RECT  1.845 1.760 2.005 2.595 ;
        RECT  1.695 1.760 1.845 1.920 ;
        RECT  1.535 0.995 1.695 1.920 ;
        RECT  1.365 2.825 1.625 3.220 ;
        RECT  1.510 0.995 1.535 1.155 ;
        RECT  1.250 0.555 1.510 1.155 ;
        RECT  0.745 2.825 1.365 2.985 ;
        RECT  0.485 2.725 0.745 2.985 ;
    END
END AOI32X4

MACRO AOI32X2
    CLASS CORE ;
    FOREIGN AOI32X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.895 1.925 4.935 2.585 ;
        RECT  4.865 0.610 4.895 2.585 ;
        RECT  4.735 0.610 4.865 2.725 ;
        RECT  3.955 0.610 4.735 0.770 ;
        RECT  4.725 1.990 4.735 2.725 ;
        RECT  4.605 2.125 4.725 2.725 ;
        RECT  3.815 2.170 4.605 2.330 ;
        RECT  3.530 0.510 3.955 0.770 ;
        RECT  3.555 2.170 3.815 2.770 ;
        RECT  1.990 0.610 3.530 0.770 ;
        RECT  1.565 0.510 1.990 0.770 ;
        END
        ANTENNADIFFAREA     1.3910 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.395 0.950 4.555 1.405 ;
        RECT  3.555 0.950 4.395 1.110 ;
        RECT  3.475 0.950 3.555 1.765 ;
        RECT  3.395 0.950 3.475 2.000 ;
        RECT  3.345 1.290 3.395 2.000 ;
        RECT  3.315 1.355 3.345 2.000 ;
        RECT  3.215 1.740 3.315 2.000 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.305 4.125 1.565 ;
        RECT  3.805 1.305 4.015 1.990 ;
        END
        ANTENNAGATEAREA     0.3536 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.265 2.785 1.525 ;
        RECT  2.585 1.265 2.635 1.580 ;
        RECT  2.425 0.950 2.585 1.580 ;
        RECT  0.855 0.950 2.425 1.110 ;
        RECT  0.695 0.950 0.855 1.520 ;
        RECT  0.625 1.360 0.695 1.520 ;
        RECT  0.365 1.360 0.625 1.665 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.795 2.475 1.955 ;
        RECT  1.105 1.700 1.255 1.990 ;
        RECT  1.045 1.700 1.105 2.005 ;
        RECT  0.845 1.745 1.045 2.005 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.290 2.010 1.580 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 -0.250 5.060 0.250 ;
        RECT  4.545 -0.250 4.805 0.405 ;
        RECT  2.985 -0.250 4.545 0.250 ;
        RECT  2.725 -0.250 2.985 0.405 ;
        RECT  0.455 -0.250 2.725 0.250 ;
        RECT  0.195 -0.250 0.455 0.935 ;
        RECT  0.000 -0.250 0.195 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.795 3.440 5.060 3.940 ;
        RECT  2.535 2.655 2.795 3.940 ;
        RECT  1.810 3.440 2.535 3.940 ;
        RECT  1.550 3.285 1.810 3.940 ;
        RECT  0.785 3.440 1.550 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.065 2.515 4.325 3.115 ;
        RECT  3.305 2.955 4.065 3.115 ;
        RECT  3.145 2.220 3.305 3.115 ;
        RECT  3.045 2.220 3.145 2.820 ;
        RECT  2.285 2.220 3.045 2.380 ;
        RECT  2.025 2.220 2.285 2.820 ;
        RECT  1.335 2.220 2.025 2.380 ;
        RECT  1.075 2.220 1.335 2.820 ;
        RECT  0.385 2.220 1.075 2.380 ;
        RECT  0.125 2.220 0.385 2.820 ;
    END
END AOI32X2

MACRO AOI32X1
    CLASS CORE ;
    FOREIGN AOI32X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.070 1.290 3.095 1.765 ;
        RECT  3.045 1.195 3.070 1.765 ;
        RECT  2.885 1.195 3.045 2.330 ;
        RECT  1.885 1.195 2.885 1.355 ;
        RECT  2.425 2.170 2.885 2.330 ;
        RECT  2.165 2.170 2.425 2.770 ;
        RECT  1.625 0.695 1.885 1.355 ;
        END
        ANTENNADIFFAREA     0.7073 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 1.550 2.695 1.990 ;
        RECT  2.355 1.550 2.400 1.810 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 1.550 2.175 1.990 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.510 1.065 1.770 ;
        RECT  0.585 1.510 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 1.550 1.545 1.810 ;
        RECT  1.285 1.010 1.445 1.810 ;
        RECT  1.255 1.010 1.285 1.170 ;
        RECT  1.045 0.880 1.255 1.170 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 -0.250 3.220 0.250 ;
        RECT  2.555 -0.250 2.815 1.015 ;
        RECT  0.385 -0.250 2.555 0.250 ;
        RECT  0.125 -0.250 0.385 1.265 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 3.440 3.220 3.940 ;
        RECT  1.145 2.510 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.170 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.835 2.510 2.935 2.770 ;
        RECT  2.675 2.510 2.835 3.110 ;
        RECT  1.915 2.950 2.675 3.110 ;
        RECT  1.755 2.170 1.915 3.110 ;
        RECT  1.655 2.170 1.755 2.770 ;
        RECT  0.895 2.170 1.655 2.330 ;
        RECT  0.635 2.170 0.895 2.770 ;
    END
END AOI32X1

MACRO AOI32XL
    CLASS CORE ;
    FOREIGN AOI32XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.070 1.290 3.095 1.765 ;
        RECT  3.045 1.210 3.070 1.765 ;
        RECT  2.885 1.210 3.045 2.330 ;
        RECT  1.915 1.210 2.885 1.370 ;
        RECT  2.425 2.170 2.885 2.330 ;
        RECT  2.265 2.170 2.425 2.705 ;
        RECT  2.165 2.445 2.265 2.705 ;
        RECT  1.755 0.780 1.915 1.370 ;
        RECT  1.655 0.780 1.755 1.040 ;
        END
        ANTENNADIFFAREA     0.3592 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.375 1.550 2.670 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 1.550 2.175 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.590 1.145 1.850 ;
        RECT  0.585 1.590 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.525 1.550 1.625 1.810 ;
        RECT  1.365 1.220 1.525 1.810 ;
        RECT  1.255 1.220 1.365 1.380 ;
        RECT  1.095 0.880 1.255 1.380 ;
        RECT  1.045 0.880 1.095 1.170 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.805 -0.250 3.220 0.250 ;
        RECT  2.545 -0.250 2.805 1.030 ;
        RECT  0.665 -0.250 2.545 0.250 ;
        RECT  0.405 -0.250 0.665 1.030 ;
        RECT  0.000 -0.250 0.405 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 3.440 3.220 3.940 ;
        RECT  1.145 2.510 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.510 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.835 2.510 2.935 2.770 ;
        RECT  2.675 2.510 2.835 3.045 ;
        RECT  1.915 2.885 2.675 3.045 ;
        RECT  1.815 2.435 1.915 3.045 ;
        RECT  1.755 2.170 1.815 3.045 ;
        RECT  1.655 2.170 1.755 2.695 ;
        RECT  0.895 2.170 1.655 2.330 ;
        RECT  0.735 2.170 0.895 2.695 ;
        RECT  0.635 2.435 0.735 2.695 ;
    END
END AOI32XL

MACRO AOI31X4
    CLASS CORE ;
    FOREIGN AOI31X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.225 4.475 2.145 ;
        RECT  4.015 1.225 4.265 1.425 ;
        RECT  4.015 1.945 4.265 2.145 ;
        RECT  3.765 0.590 4.015 1.425 ;
        RECT  3.965 1.945 4.015 2.585 ;
        RECT  3.705 1.945 3.965 3.080 ;
        RECT  3.705 0.590 3.765 1.190 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 1.440 2.175 1.990 ;
        END
        ANTENNAGATEAREA     0.0975 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.475 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.825 1.510 1.075 1.770 ;
        RECT  0.585 1.510 0.825 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 1.700 1.715 1.990 ;
        RECT  1.295 1.510 1.555 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 -0.250 4.600 0.250 ;
        RECT  4.215 -0.250 4.475 1.045 ;
        RECT  3.455 -0.250 4.215 0.250 ;
        RECT  3.195 -0.250 3.455 1.095 ;
        RECT  2.305 -0.250 3.195 0.250 ;
        RECT  2.045 -0.250 2.305 0.850 ;
        RECT  0.385 -0.250 2.045 0.250 ;
        RECT  0.125 -0.250 0.385 1.165 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 3.440 4.600 3.940 ;
        RECT  4.215 2.325 4.475 3.940 ;
        RECT  3.455 3.440 4.215 3.940 ;
        RECT  3.195 2.275 3.455 3.940 ;
        RECT  1.305 3.440 3.195 3.940 ;
        RECT  1.045 2.835 1.305 3.940 ;
        RECT  0.385 3.440 1.045 3.940 ;
        RECT  0.125 2.835 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.975 1.605 4.085 1.765 ;
        RECT  2.895 1.150 2.975 2.160 ;
        RECT  2.815 0.695 2.895 3.205 ;
        RECT  2.735 0.695 2.815 1.310 ;
        RECT  2.735 2.000 2.815 3.205 ;
        RECT  2.515 1.510 2.635 1.770 ;
        RECT  2.355 1.100 2.515 2.330 ;
        RECT  1.725 1.100 2.355 1.260 ;
        RECT  2.335 2.170 2.355 2.330 ;
        RECT  2.075 2.170 2.335 2.430 ;
        RECT  1.565 2.170 1.825 2.430 ;
        RECT  1.465 1.000 1.725 1.260 ;
        RECT  0.785 2.170 1.565 2.330 ;
        RECT  0.525 2.170 0.785 2.430 ;
    END
END AOI31X4

MACRO AOI31X2
    CLASS CORE ;
    FOREIGN AOI31X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 1.515 4.015 2.175 ;
        RECT  3.805 1.130 3.965 2.750 ;
        RECT  3.245 1.130 3.805 1.290 ;
        RECT  3.695 2.490 3.805 2.750 ;
        RECT  2.985 0.690 3.245 1.290 ;
        RECT  0.610 0.950 2.985 1.110 ;
        RECT  0.605 0.690 0.610 1.110 ;
        RECT  0.345 0.690 0.605 1.290 ;
        END
        ANTENNADIFFAREA     0.9414 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.325 1.510 3.585 2.120 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.400 2.045 1.660 ;
        RECT  1.505 1.290 1.715 1.660 ;
        RECT  1.445 1.400 1.505 1.660 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.305 1.740 2.565 2.000 ;
        RECT  1.255 1.840 2.305 2.000 ;
        RECT  1.045 1.290 1.255 2.000 ;
        RECT  0.895 1.740 1.045 2.000 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 1.680 3.105 1.940 ;
        RECT  3.005 1.680 3.095 1.990 ;
        RECT  2.845 1.680 3.005 2.340 ;
        RECT  0.555 2.180 2.845 2.340 ;
        RECT  0.395 1.725 0.555 2.340 ;
        RECT  0.335 1.725 0.395 1.990 ;
        RECT  0.295 1.725 0.335 1.985 ;
        END
        ANTENNAGATEAREA     0.3900 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.785 -0.250 4.600 0.250 ;
        RECT  3.525 -0.250 3.785 0.945 ;
        RECT  1.905 -0.250 3.525 0.250 ;
        RECT  1.645 -0.250 1.905 0.765 ;
        RECT  0.000 -0.250 1.645 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 3.440 4.600 3.940 ;
        RECT  2.675 2.860 2.935 3.940 ;
        RECT  1.915 3.440 2.675 3.940 ;
        RECT  1.655 2.860 1.915 3.940 ;
        RECT  0.895 3.440 1.655 3.940 ;
        RECT  0.635 2.860 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.205 2.420 4.465 3.090 ;
        RECT  3.445 2.930 4.205 3.090 ;
        RECT  3.185 2.420 3.445 3.090 ;
        RECT  2.425 2.520 3.185 2.680 ;
        RECT  2.165 2.520 2.425 3.120 ;
        RECT  1.405 2.520 2.165 2.680 ;
        RECT  1.145 2.520 1.405 3.120 ;
        RECT  0.385 2.520 1.145 2.680 ;
        RECT  0.125 2.520 0.385 3.120 ;
    END
END AOI31X2

MACRO AOI31X1
    CLASS CORE ;
    FOREIGN AOI31X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.350 2.635 2.400 ;
        RECT  2.425 1.110 2.560 2.475 ;
        RECT  2.400 1.110 2.425 2.915 ;
        RECT  1.710 1.110 2.400 1.270 ;
        RECT  2.165 2.315 2.400 2.915 ;
        RECT  1.450 1.010 1.710 1.270 ;
        END
        ANTENNADIFFAREA     0.5594 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 1.510 2.215 1.990 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.820 1.760 1.065 2.020 ;
        RECT  0.805 1.500 0.820 2.020 ;
        RECT  0.585 1.500 0.805 1.990 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 1.450 1.715 1.990 ;
        RECT  1.315 1.450 1.465 1.710 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 -0.250 2.760 0.250 ;
        RECT  2.225 -0.250 2.485 0.870 ;
        RECT  0.510 -0.250 2.225 0.250 ;
        RECT  0.250 -0.250 0.510 1.265 ;
        RECT  0.000 -0.250 0.250 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 3.440 2.760 3.940 ;
        RECT  1.145 2.585 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.415 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.655 2.205 1.915 2.915 ;
        RECT  0.895 2.205 1.655 2.365 ;
        RECT  0.635 2.205 0.895 2.915 ;
    END
END AOI31X1

MACRO AOI31XL
    CLASS CORE ;
    FOREIGN AOI31XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.515 1.515 2.635 2.400 ;
        RECT  2.425 1.130 2.515 2.625 ;
        RECT  2.355 1.130 2.425 2.715 ;
        RECT  1.785 1.130 2.355 1.290 ;
        RECT  2.165 2.455 2.355 2.715 ;
        RECT  1.525 1.030 1.785 1.290 ;
        END
        ANTENNADIFFAREA     0.3160 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 1.510 2.175 1.990 ;
        END
        ANTENNAGATEAREA     0.0871 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.805 1.725 1.065 1.985 ;
        RECT  0.585 1.510 0.805 1.990 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.510 1.715 1.990 ;
        RECT  1.285 1.510 1.505 1.770 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 -0.250 2.760 0.250 ;
        RECT  2.095 -0.250 2.355 0.870 ;
        RECT  0.580 -0.250 2.095 0.250 ;
        RECT  0.320 -0.250 0.580 1.230 ;
        RECT  0.000 -0.250 0.320 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 3.440 2.760 3.940 ;
        RECT  1.145 2.515 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.435 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.815 2.455 1.915 2.715 ;
        RECT  1.655 2.175 1.815 2.715 ;
        RECT  0.895 2.175 1.655 2.335 ;
        RECT  0.735 2.175 0.895 2.715 ;
        RECT  0.635 2.455 0.735 2.715 ;
    END
END AOI31XL

MACRO AOI222X4
    CLASS CORE ;
    FOREIGN AOI222X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.345 1.105 5.395 2.135 ;
        RECT  5.285 1.035 5.345 2.135 ;
        RECT  5.185 0.600 5.285 3.065 ;
        RECT  5.025 0.600 5.185 1.200 ;
        RECT  5.125 1.975 5.185 3.065 ;
        RECT  5.025 2.125 5.125 3.065 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.560 0.925 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.510 2.065 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.285 1.510 2.635 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.275 1.450 3.555 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 1.450 3.095 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.835 -0.250 5.980 0.250 ;
        RECT  5.575 -0.250 5.835 1.185 ;
        RECT  4.775 -0.250 5.575 0.250 ;
        RECT  4.515 -0.250 4.775 1.095 ;
        RECT  3.755 -0.250 4.515 0.250 ;
        RECT  3.495 -0.250 3.755 0.825 ;
        RECT  1.590 -0.250 3.495 0.250 ;
        RECT  1.330 -0.250 1.590 0.825 ;
        RECT  0.000 -0.250 1.330 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.795 3.440 5.980 3.940 ;
        RECT  5.535 2.275 5.795 3.940 ;
        RECT  4.775 3.440 5.535 3.940 ;
        RECT  4.515 2.615 4.775 3.940 ;
        RECT  1.185 3.440 4.515 3.940 ;
        RECT  0.925 3.285 1.185 3.940 ;
        RECT  0.385 3.440 0.925 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.825 1.510 4.925 1.770 ;
        RECT  4.665 1.275 4.825 2.435 ;
        RECT  4.265 1.275 4.665 1.435 ;
        RECT  4.265 2.275 4.665 2.435 ;
        RECT  3.895 1.650 4.435 1.910 ;
        RECT  4.105 0.655 4.265 1.435 ;
        RECT  4.105 2.275 4.265 3.110 ;
        RECT  4.005 0.655 4.105 0.915 ;
        RECT  4.005 2.510 4.105 3.110 ;
        RECT  3.735 1.095 3.895 2.330 ;
        RECT  2.770 1.095 3.735 1.255 ;
        RECT  3.225 2.170 3.735 2.330 ;
        RECT  3.475 2.510 3.735 2.770 ;
        RECT  2.715 2.610 3.475 2.770 ;
        RECT  2.965 2.170 3.225 2.430 ;
        RECT  2.510 0.995 2.770 1.255 ;
        RECT  2.455 2.170 2.715 2.770 ;
        RECT  0.475 1.095 2.510 1.255 ;
        RECT  1.695 2.610 2.455 2.770 ;
        RECT  1.945 2.170 2.205 2.430 ;
        RECT  0.785 2.170 1.945 2.330 ;
        RECT  1.435 2.510 1.695 2.770 ;
        RECT  0.525 2.170 0.785 2.770 ;
        RECT  0.215 0.995 0.475 1.255 ;
    END
END AOI222X4

MACRO AOI222X2
    CLASS CORE ;
    FOREIGN AOI222X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 0.945 7.235 1.990 ;
        RECT  7.025 0.945 7.185 2.260 ;
        RECT  6.130 0.945 7.025 1.105 ;
        RECT  6.505 2.100 7.025 2.260 ;
        RECT  6.245 2.100 6.505 2.700 ;
        RECT  5.485 2.100 6.245 2.260 ;
        RECT  5.735 0.840 6.130 1.105 ;
        RECT  3.955 0.945 5.735 1.105 ;
        RECT  5.225 2.100 5.485 2.700 ;
        RECT  3.530 0.845 3.955 1.105 ;
        RECT  1.530 0.945 3.530 1.105 ;
        RECT  1.145 0.845 1.530 1.105 ;
        END
        ANTENNADIFFAREA     1.4954 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.055 1.290 2.175 1.580 ;
        RECT  1.965 1.290 2.055 1.650 ;
        RECT  1.795 1.310 1.965 1.650 ;
        RECT  0.755 1.310 1.795 1.470 ;
        RECT  0.595 1.310 0.755 1.770 ;
        RECT  0.495 1.510 0.595 1.770 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.650 1.575 1.810 ;
        RECT  1.045 1.650 1.255 1.990 ;
        RECT  0.975 1.650 1.045 1.810 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.535 1.510 4.635 1.770 ;
        RECT  4.375 1.510 4.535 1.920 ;
        RECT  3.095 1.760 4.375 1.920 ;
        RECT  2.935 1.290 3.095 1.920 ;
        RECT  2.885 1.290 2.935 1.770 ;
        RECT  2.835 1.510 2.885 1.770 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.320 4.125 1.580 ;
        RECT  3.805 1.290 4.015 1.580 ;
        RECT  3.525 1.320 3.805 1.580 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.415 1.510 6.675 1.920 ;
        RECT  5.395 1.760 6.415 1.920 ;
        RECT  5.235 1.290 5.395 1.920 ;
        RECT  5.185 1.290 5.235 1.770 ;
        RECT  5.085 1.510 5.185 1.770 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.320 6.175 1.580 ;
        RECT  5.645 1.290 5.855 1.580 ;
        RECT  5.575 1.320 5.645 1.580 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 -0.250 7.360 0.250 ;
        RECT  6.600 -0.250 6.860 0.745 ;
        RECT  4.975 -0.250 6.600 0.250 ;
        RECT  4.715 -0.250 4.975 0.745 ;
        RECT  3.035 -0.250 4.715 0.250 ;
        RECT  2.775 -0.250 3.035 0.745 ;
        RECT  2.325 -0.250 2.775 0.250 ;
        RECT  2.065 -0.250 2.325 0.745 ;
        RECT  0.485 -0.250 2.065 0.250 ;
        RECT  0.225 -0.250 0.485 1.130 ;
        RECT  0.000 -0.250 0.225 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 3.440 7.360 3.940 ;
        RECT  2.165 2.465 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.755 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.080 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.755 2.465 7.015 3.040 ;
        RECT  5.995 2.880 6.755 3.040 ;
        RECT  5.735 2.465 5.995 3.040 ;
        RECT  4.975 2.880 5.735 3.040 ;
        RECT  4.715 2.080 4.975 3.040 ;
        RECT  3.955 2.880 4.715 3.040 ;
        RECT  4.205 2.100 4.465 2.700 ;
        RECT  3.445 2.100 4.205 2.260 ;
        RECT  3.695 2.465 3.955 3.040 ;
        RECT  2.935 2.880 3.695 3.040 ;
        RECT  3.185 2.100 3.445 2.700 ;
        RECT  1.915 2.100 3.185 2.260 ;
        RECT  2.675 2.465 2.935 3.040 ;
        RECT  1.655 2.080 1.915 3.020 ;
        RECT  0.895 2.170 1.655 2.330 ;
        RECT  0.635 2.170 0.895 2.770 ;
    END
END AOI222X2

MACRO AOI222X1
    CLASS CORE ;
    FOREIGN AOI222X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 0.950 4.015 1.990 ;
        RECT  3.805 0.950 3.990 2.130 ;
        RECT  2.910 0.950 3.805 1.110 ;
        RECT  3.445 1.970 3.805 2.130 ;
        RECT  3.285 1.970 3.445 2.740 ;
        RECT  3.185 2.140 3.285 2.740 ;
        RECT  2.585 0.850 2.910 1.110 ;
        RECT  0.610 0.950 2.585 1.110 ;
        RECT  0.325 0.850 0.610 1.110 ;
        END
        ANTENNADIFFAREA     0.9478 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.040 1.290 1.300 1.770 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.295 1.290 0.555 1.750 ;
        RECT  0.125 1.290 0.295 1.580 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.290 1.785 1.770 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.290 2.595 1.770 ;
        RECT  1.965 1.290 2.335 1.580 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.320 1.290 3.615 1.790 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 1.290 3.095 1.770 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.785 -0.250 4.140 0.250 ;
        RECT  3.525 -0.250 3.785 0.770 ;
        RECT  1.665 -0.250 3.525 0.250 ;
        RECT  1.405 -0.250 1.665 0.745 ;
        RECT  0.000 -0.250 1.405 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 3.440 4.140 3.940 ;
        RECT  1.145 2.420 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.080 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.695 2.420 3.955 3.090 ;
        RECT  2.935 2.930 3.695 3.090 ;
        RECT  2.675 2.080 2.935 3.090 ;
        RECT  1.915 2.930 2.675 3.090 ;
        RECT  2.325 2.140 2.425 2.740 ;
        RECT  2.165 1.970 2.325 2.740 ;
        RECT  0.895 1.970 2.165 2.130 ;
        RECT  1.655 2.420 1.915 3.090 ;
        RECT  0.635 1.970 0.895 3.020 ;
    END
END AOI222X1

MACRO AOI222XL
    CLASS CORE ;
    FOREIGN AOI222XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.415 0.925 3.575 2.440 ;
        RECT  2.545 0.925 3.415 1.085 ;
        RECT  3.345 1.700 3.415 2.440 ;
        RECT  3.155 2.280 3.345 2.440 ;
        RECT  2.895 2.280 3.155 2.540 ;
        RECT  2.285 0.820 2.545 1.085 ;
        RECT  0.610 0.925 2.285 1.085 ;
        RECT  0.325 0.820 0.610 1.085 ;
        END
        ANTENNADIFFAREA     0.4653 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.865 1.850 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.405 1.770 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.525 1.510 1.785 1.770 ;
        RECT  1.255 1.510 1.525 1.670 ;
        RECT  1.045 1.290 1.255 1.670 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.245 1.265 2.345 1.525 ;
        RECT  1.965 1.265 2.245 1.840 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.145 1.265 3.235 1.455 ;
        RECT  2.815 1.265 3.145 1.585 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.775 2.915 2.055 ;
        RECT  2.425 1.700 2.635 2.055 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.505 -0.250 3.680 0.250 ;
        RECT  3.245 -0.250 3.505 0.745 ;
        RECT  1.505 -0.250 3.245 0.250 ;
        RECT  1.245 -0.250 1.505 0.745 ;
        RECT  0.000 -0.250 1.245 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 3.440 3.680 3.940 ;
        RECT  0.925 3.285 1.185 3.940 ;
        RECT  0.385 3.440 0.925 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.295 2.955 3.555 3.215 ;
        RECT  2.670 2.955 3.295 3.115 ;
        RECT  2.410 2.955 2.670 3.215 ;
        RECT  1.695 2.955 2.410 3.115 ;
        RECT  1.945 2.035 2.205 2.360 ;
        RECT  0.785 2.035 1.945 2.195 ;
        RECT  1.535 2.375 1.695 3.115 ;
        RECT  1.435 2.375 1.535 2.635 ;
        RECT  0.625 2.035 0.785 2.680 ;
        RECT  0.525 2.420 0.625 2.680 ;
    END
END AOI222XL

MACRO AOI221X4
    CLASS CORE ;
    FOREIGN AOI221X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.345 1.255 5.395 2.175 ;
        RECT  5.185 1.255 5.345 2.370 ;
        RECT  4.755 1.255 5.185 1.415 ;
        RECT  4.755 2.210 5.185 2.370 ;
        RECT  4.495 0.675 4.755 1.415 ;
        RECT  4.495 2.210 4.755 3.150 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.560 2.885 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.610 0.925 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.415 2.245 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 1.530 1.765 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.265 -0.250 5.520 0.250 ;
        RECT  5.005 -0.250 5.265 1.075 ;
        RECT  4.245 -0.250 5.005 0.250 ;
        RECT  3.985 -0.250 4.245 0.815 ;
        RECT  2.650 -0.250 3.985 0.250 ;
        RECT  2.390 -0.250 2.650 0.805 ;
        RECT  0.775 -0.250 2.390 0.250 ;
        RECT  0.515 -0.250 0.775 1.255 ;
        RECT  0.000 -0.250 0.515 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.265 3.440 5.520 3.940 ;
        RECT  5.005 2.615 5.265 3.940 ;
        RECT  4.245 3.440 5.005 3.940 ;
        RECT  3.985 2.325 4.245 3.940 ;
        RECT  1.185 3.440 3.985 3.940 ;
        RECT  0.925 3.285 1.185 3.940 ;
        RECT  0.385 3.440 0.925 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.245 1.605 4.925 1.865 ;
        RECT  4.085 1.005 4.245 2.145 ;
        RECT  3.735 1.005 4.085 1.165 ;
        RECT  3.735 1.985 4.085 2.145 ;
        RECT  3.645 1.545 3.905 1.805 ;
        RECT  3.475 0.565 3.735 1.165 ;
        RECT  3.475 1.985 3.735 2.925 ;
        RECT  3.225 1.595 3.645 1.755 ;
        RECT  3.065 1.035 3.225 2.760 ;
        RECT  2.965 1.035 3.065 1.295 ;
        RECT  2.965 2.160 3.065 2.760 ;
        RECT  1.595 1.065 2.965 1.225 ;
        RECT  2.615 2.170 2.715 2.770 ;
        RECT  2.455 2.170 2.615 3.110 ;
        RECT  1.695 2.950 2.455 3.110 ;
        RECT  1.945 2.170 2.205 2.770 ;
        RECT  0.785 2.170 1.945 2.330 ;
        RECT  1.535 2.510 1.695 3.110 ;
        RECT  1.335 1.010 1.595 1.270 ;
        RECT  1.435 2.510 1.535 2.770 ;
        RECT  0.625 2.170 0.785 2.545 ;
        RECT  0.525 2.285 0.625 2.545 ;
    END
END AOI221X4

MACRO AOI221X2
    CLASS CORE ;
    FOREIGN AOI221X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 2.170 5.305 2.770 ;
        RECT  5.045 1.740 5.205 2.770 ;
        RECT  4.935 0.910 5.165 1.170 ;
        RECT  4.935 1.740 5.045 1.900 ;
        RECT  4.905 0.910 4.935 1.900 ;
        RECT  4.775 0.950 4.905 1.900 ;
        RECT  3.645 0.950 4.775 1.110 ;
        RECT  4.725 1.290 4.775 1.580 ;
        RECT  3.385 0.850 3.645 1.110 ;
        RECT  2.255 0.950 3.385 1.110 ;
        RECT  2.095 0.755 2.255 1.110 ;
        RECT  1.475 0.755 2.095 0.915 ;
        RECT  1.215 0.655 1.475 0.915 ;
        END
        ANTENNADIFFAREA     1.1712 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.385 1.290 5.855 1.715 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 1.290 2.175 1.580 ;
        RECT  1.915 1.290 2.125 1.680 ;
        RECT  1.865 1.095 1.915 1.680 ;
        RECT  1.755 1.095 1.865 1.450 ;
        RECT  0.795 1.095 1.755 1.255 ;
        RECT  0.725 1.095 0.795 1.765 ;
        RECT  0.565 1.095 0.725 1.905 ;
        RECT  0.465 1.515 0.565 1.905 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.440 1.575 1.700 ;
        RECT  1.045 1.440 1.255 1.990 ;
        RECT  0.975 1.440 1.045 1.700 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.325 1.515 4.425 1.790 ;
        RECT  4.165 1.290 4.325 1.790 ;
        RECT  3.095 1.290 4.165 1.450 ;
        RECT  2.925 1.290 3.095 1.580 ;
        RECT  2.665 1.290 2.925 1.680 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.650 3.945 1.810 ;
        RECT  3.345 1.650 3.555 1.990 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.675 -0.250 5.980 0.250 ;
        RECT  5.415 -0.250 5.675 1.110 ;
        RECT  4.625 -0.250 5.415 0.250 ;
        RECT  4.365 -0.250 4.625 0.770 ;
        RECT  2.695 -0.250 4.365 0.250 ;
        RECT  2.435 -0.250 2.695 0.770 ;
        RECT  0.585 -0.250 2.435 0.250 ;
        RECT  0.325 -0.250 0.585 0.915 ;
        RECT  0.000 -0.250 0.325 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 3.440 5.980 3.940 ;
        RECT  2.095 2.955 2.355 3.940 ;
        RECT  1.435 3.440 2.095 3.940 ;
        RECT  1.175 3.285 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.255 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.555 2.080 5.815 3.110 ;
        RECT  4.795 2.950 5.555 3.110 ;
        RECT  4.535 2.080 4.795 3.110 ;
        RECT  3.775 2.950 4.535 3.110 ;
        RECT  4.025 2.170 4.285 2.770 ;
        RECT  3.265 2.170 4.025 2.330 ;
        RECT  3.515 2.510 3.775 3.110 ;
        RECT  2.755 2.950 3.515 3.110 ;
        RECT  3.165 2.170 3.265 2.770 ;
        RECT  3.005 2.105 3.165 2.770 ;
        RECT  1.835 2.105 3.005 2.265 ;
        RECT  2.595 2.445 2.755 3.110 ;
        RECT  2.495 2.445 2.595 2.705 ;
        RECT  1.675 2.105 1.835 2.820 ;
        RECT  1.575 2.220 1.675 2.820 ;
        RECT  0.895 2.220 1.575 2.380 ;
        RECT  0.635 2.220 0.895 3.160 ;
    END
END AOI221X2

MACRO AOI221X1
    CLASS CORE ;
    FOREIGN AOI221X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.475 1.105 3.555 2.585 ;
        RECT  3.315 0.850 3.475 3.020 ;
        RECT  3.215 0.850 3.315 1.110 ;
        RECT  3.215 2.080 3.315 3.020 ;
        RECT  1.990 0.950 3.215 1.110 ;
        RECT  1.715 0.850 1.990 1.110 ;
        END
        ANTENNADIFFAREA     0.7686 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.875 1.290 3.135 1.860 ;
        END
        ANTENNAGATEAREA     0.1963 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.515 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.700 1.035 1.985 ;
        RECT  0.585 1.700 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.365 1.290 2.635 1.765 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.420 2.145 1.680 ;
        RECT  1.510 1.290 1.715 1.680 ;
        RECT  1.505 1.290 1.510 1.580 ;
        END
        ANTENNAGATEAREA     0.2171 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.915 -0.250 3.680 0.250 ;
        RECT  2.655 -0.250 2.915 0.770 ;
        RECT  1.095 -0.250 2.655 0.250 ;
        RECT  0.835 -0.250 1.095 1.110 ;
        RECT  0.000 -0.250 0.835 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 3.440 3.680 3.940 ;
        RECT  1.175 2.555 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.255 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.705 2.080 2.965 3.020 ;
        RECT  1.945 2.860 2.705 3.020 ;
        RECT  2.195 2.075 2.455 2.675 ;
        RECT  1.410 2.075 2.195 2.235 ;
        RECT  1.685 2.420 1.945 3.020 ;
        RECT  1.250 2.075 1.410 2.375 ;
        RECT  0.895 2.215 1.250 2.375 ;
        RECT  0.635 2.215 0.895 3.195 ;
    END
END AOI221X1

MACRO AOI221XL
    CLASS CORE ;
    FOREIGN AOI221XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.045 1.105 3.095 2.175 ;
        RECT  2.885 0.850 3.045 2.475 ;
        RECT  2.700 0.850 2.885 1.110 ;
        RECT  2.785 2.215 2.885 2.475 ;
        RECT  1.530 0.950 2.700 1.110 ;
        RECT  1.145 0.850 1.530 1.110 ;
        END
        ANTENNADIFFAREA     0.4234 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.330 2.670 1.590 ;
        RECT  2.595 1.290 2.635 1.765 ;
        RECT  2.425 1.290 2.595 1.955 ;
        RECT  2.410 1.330 2.425 1.955 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.515 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.875 0.875 2.165 ;
        RECT  0.585 1.625 0.795 2.165 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.065 1.290 2.175 1.580 ;
        RECT  1.795 1.290 2.065 1.765 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 1.420 1.575 1.680 ;
        RECT  1.255 1.420 1.315 1.580 ;
        RECT  1.045 1.290 1.255 1.580 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.320 -0.250 3.220 0.250 ;
        RECT  2.060 -0.250 2.320 0.770 ;
        RECT  0.585 -0.250 2.060 0.250 ;
        RECT  0.325 -0.250 0.585 1.110 ;
        RECT  0.000 -0.250 0.325 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 3.440 3.220 3.940 ;
        RECT  0.925 3.285 1.185 3.940 ;
        RECT  0.385 3.440 0.925 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.235 2.880 2.495 3.140 ;
        RECT  1.695 2.930 2.235 3.090 ;
        RECT  1.995 2.215 2.095 2.475 ;
        RECT  1.835 2.015 1.995 2.475 ;
        RECT  1.265 2.015 1.835 2.175 ;
        RECT  1.435 2.880 1.695 3.140 ;
        RECT  1.105 2.015 1.265 2.575 ;
        RECT  0.785 2.415 1.105 2.575 ;
        RECT  0.525 2.415 0.785 2.675 ;
    END
END AOI221XL

MACRO AOI22X4
    CLASS CORE ;
    FOREIGN AOI22X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.305 1.105 6.315 1.765 ;
        RECT  6.105 1.025 6.305 2.310 ;
        RECT  5.785 1.025 6.105 1.225 ;
        RECT  5.785 2.110 6.105 2.310 ;
        RECT  5.455 0.625 5.785 1.225 ;
        RECT  5.555 2.110 5.785 2.770 ;
        RECT  5.525 2.170 5.555 2.770 ;
        RECT  4.765 2.170 5.525 2.370 ;
        RECT  5.395 0.625 5.455 1.170 ;
        RECT  5.185 0.470 5.395 1.170 ;
        RECT  4.085 0.925 5.185 1.125 ;
        RECT  4.505 2.170 4.765 2.770 ;
        RECT  3.745 2.170 4.505 2.370 ;
        RECT  3.825 0.495 4.085 1.125 ;
        RECT  2.285 0.590 3.825 0.790 ;
        RECT  3.485 2.170 3.745 2.770 ;
        RECT  2.025 0.590 2.285 0.870 ;
        RECT  0.385 0.590 2.025 0.790 ;
        RECT  0.125 0.475 0.385 1.075 ;
        END
        ANTENNADIFFAREA     2.3729 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.375 2.935 1.635 ;
        RECT  2.585 1.375 2.635 1.990 ;
        RECT  2.425 1.155 2.585 1.990 ;
        RECT  1.445 1.155 2.425 1.315 ;
        RECT  1.285 1.155 1.445 1.565 ;
        RECT  0.775 1.405 1.285 1.565 ;
        END
        ANTENNAGATEAREA     0.7254 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.495 2.245 1.755 ;
        RECT  2.145 1.495 2.150 1.765 ;
        RECT  1.985 1.495 2.145 1.905 ;
        RECT  0.555 1.745 1.985 1.905 ;
        RECT  0.395 1.515 0.555 1.905 ;
        RECT  0.335 1.515 0.395 1.775 ;
        RECT  0.295 1.290 0.335 1.775 ;
        RECT  0.125 1.290 0.295 1.770 ;
        END
        ANTENNAGATEAREA     0.7254 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.335 4.735 1.595 ;
        RECT  3.575 1.340 4.475 1.500 ;
        RECT  3.555 1.340 3.575 1.915 ;
        RECT  3.345 1.290 3.555 1.915 ;
        RECT  3.315 1.655 3.345 1.915 ;
        END
        ANTENNAGATEAREA     0.7371 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.665 1.600 5.925 1.860 ;
        RECT  5.210 1.700 5.665 1.860 ;
        RECT  4.975 1.700 5.210 1.940 ;
        RECT  4.085 1.780 4.975 1.940 ;
        RECT  4.015 1.680 4.085 1.940 ;
        RECT  3.825 1.680 4.015 1.990 ;
        RECT  3.805 1.700 3.825 1.990 ;
        END
        ANTENNAGATEAREA     0.7371 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 -0.250 6.440 0.250 ;
        RECT  4.675 -0.250 4.935 0.745 ;
        RECT  3.185 -0.250 4.675 0.250 ;
        RECT  2.925 -0.250 3.185 0.405 ;
        RECT  1.350 -0.250 2.925 0.250 ;
        RECT  1.090 -0.250 1.350 0.405 ;
        RECT  0.000 -0.250 1.090 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.685 3.440 6.440 3.940 ;
        RECT  2.425 3.285 2.685 3.940 ;
        RECT  1.885 3.440 2.425 3.940 ;
        RECT  1.625 3.285 1.885 3.940 ;
        RECT  0.935 3.440 1.625 3.940 ;
        RECT  0.675 3.285 0.935 3.940 ;
        RECT  0.000 3.440 0.675 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.035 2.490 6.295 3.110 ;
        RECT  5.275 2.950 6.035 3.110 ;
        RECT  5.015 2.610 5.275 3.110 ;
        RECT  4.255 2.950 5.015 3.110 ;
        RECT  3.995 2.610 4.255 3.110 ;
        RECT  3.235 2.950 3.995 3.110 ;
        RECT  3.075 2.170 3.235 3.110 ;
        RECT  2.975 2.170 3.075 2.770 ;
        RECT  2.285 2.170 2.975 2.330 ;
        RECT  2.025 2.170 2.285 2.770 ;
        RECT  1.335 2.170 2.025 2.330 ;
        RECT  1.075 2.085 1.335 2.685 ;
        RECT  0.385 2.085 1.075 2.245 ;
        RECT  0.125 2.085 0.385 2.685 ;
    END
END AOI22X4

MACRO AOI22X2
    CLASS CORE ;
    FOREIGN AOI22X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.275 0.930 4.435 2.015 ;
        RECT  3.245 0.930 4.275 1.090 ;
        RECT  4.015 1.855 4.275 2.015 ;
        RECT  3.955 1.855 4.015 2.400 ;
        RECT  3.805 1.855 3.955 2.770 ;
        RECT  3.695 2.170 3.805 2.770 ;
        RECT  2.935 2.170 3.695 2.330 ;
        RECT  2.985 0.830 3.245 1.090 ;
        RECT  1.345 0.930 2.985 1.090 ;
        RECT  2.675 2.170 2.935 2.770 ;
        RECT  1.085 0.830 1.345 1.090 ;
        END
        ANTENNADIFFAREA     1.1140 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 1.510 2.055 1.770 ;
        RECT  1.795 1.270 1.955 1.770 ;
        RECT  0.695 1.270 1.795 1.430 ;
        RECT  0.535 1.270 0.695 1.770 ;
        RECT  0.435 1.510 0.535 1.770 ;
        RECT  0.335 1.610 0.435 1.770 ;
        RECT  0.125 1.610 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.610 1.515 1.870 ;
        RECT  1.045 1.610 1.255 1.990 ;
        RECT  0.915 1.610 1.045 1.870 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.995 1.415 4.095 1.675 ;
        RECT  3.835 1.270 3.995 1.675 ;
        RECT  2.635 1.270 3.835 1.430 ;
        RECT  2.475 1.270 2.635 1.990 ;
        RECT  2.425 1.510 2.475 1.990 ;
        RECT  2.335 1.510 2.425 1.770 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 1.610 3.325 1.990 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.165 -0.250 4.600 0.250 ;
        RECT  3.905 -0.250 4.165 0.745 ;
        RECT  2.325 -0.250 3.905 0.250 ;
        RECT  2.065 -0.250 2.325 0.745 ;
        RECT  0.525 -0.250 2.065 0.250 ;
        RECT  0.265 -0.250 0.525 1.015 ;
        RECT  0.000 -0.250 0.265 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 3.440 4.600 3.940 ;
        RECT  1.655 2.510 1.915 3.940 ;
        RECT  0.895 3.440 1.655 3.940 ;
        RECT  0.635 2.510 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.365 2.195 4.465 2.780 ;
        RECT  4.205 2.195 4.365 3.110 ;
        RECT  3.445 2.950 4.205 3.110 ;
        RECT  3.185 2.510 3.445 3.110 ;
        RECT  2.425 2.950 3.185 3.110 ;
        RECT  2.265 2.170 2.425 3.110 ;
        RECT  2.165 2.170 2.265 2.770 ;
        RECT  1.405 2.170 2.165 2.330 ;
        RECT  1.145 2.170 1.405 2.770 ;
        RECT  0.385 2.170 1.145 2.330 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END AOI22X2

MACRO AOI22X1
    CLASS CORE ;
    FOREIGN AOI22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.515 2.635 2.175 ;
        RECT  2.425 1.345 2.585 2.380 ;
        RECT  1.305 1.345 2.425 1.505 ;
        RECT  1.915 2.220 2.425 2.380 ;
        RECT  1.655 2.220 1.915 2.820 ;
        RECT  1.145 0.895 1.305 1.505 ;
        RECT  0.975 0.895 1.145 1.155 ;
        END
        ANTENNADIFFAREA     0.5744 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.115 1.460 0.375 1.990 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.700 1.035 1.990 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 1.690 2.245 2.040 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.285 1.700 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.255 -0.250 2.760 0.250 ;
        RECT  1.995 -0.250 2.255 1.165 ;
        RECT  0.385 -0.250 1.995 0.250 ;
        RECT  0.125 -0.250 0.385 1.155 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 3.440 2.760 3.940 ;
        RECT  0.635 2.710 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.325 2.710 2.425 2.970 ;
        RECT  2.165 2.710 2.325 3.160 ;
        RECT  1.405 3.000 2.165 3.160 ;
        RECT  1.245 2.170 1.405 3.160 ;
        RECT  1.145 2.170 1.245 2.770 ;
        RECT  0.385 2.170 1.145 2.330 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END AOI22X1

MACRO AOI22XL
    CLASS CORE ;
    FOREIGN AOI22XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.515 2.635 1.990 ;
        RECT  2.425 1.010 2.585 2.330 ;
        RECT  1.235 1.010 2.425 1.170 ;
        RECT  1.915 2.170 2.425 2.330 ;
        RECT  1.755 2.170 1.915 2.630 ;
        RECT  1.655 2.370 1.755 2.630 ;
        RECT  0.975 0.910 1.235 1.170 ;
        END
        ANTENNADIFFAREA     0.3074 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.120 1.460 0.395 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.700 1.035 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 1.445 2.185 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.285 1.700 1.715 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.255 -0.250 2.760 0.250 ;
        RECT  1.995 -0.250 2.255 0.830 ;
        RECT  0.385 -0.250 1.995 0.250 ;
        RECT  0.125 -0.250 0.385 1.170 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 3.440 2.760 3.940 ;
        RECT  0.635 2.510 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.325 2.515 2.425 2.775 ;
        RECT  2.165 2.515 2.325 2.970 ;
        RECT  1.405 2.810 2.165 2.970 ;
        RECT  1.305 2.440 1.405 2.970 ;
        RECT  1.245 2.170 1.305 2.970 ;
        RECT  1.145 2.170 1.245 2.700 ;
        RECT  0.385 2.170 1.145 2.330 ;
        RECT  0.225 2.170 0.385 2.700 ;
        RECT  0.125 2.440 0.225 2.700 ;
    END
END AOI22XL

MACRO AOI211X4
    CLASS CORE ;
    FOREIGN AOI211X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.755 0.935 4.015 2.230 ;
        RECT  3.555 0.935 3.755 1.195 ;
        RECT  3.555 1.970 3.755 2.230 ;
        RECT  3.505 0.695 3.555 1.195 ;
        RECT  3.505 1.970 3.555 2.585 ;
        RECT  3.245 0.545 3.505 1.195 ;
        RECT  3.245 1.970 3.505 2.915 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 1.535 1.475 1.990 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 2.930 2.175 3.220 ;
        RECT  1.640 2.750 1.985 3.220 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.510 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 0.470 1.045 0.850 ;
        END
        ANTENNAGATEAREA     0.1287 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 -0.250 4.140 0.250 ;
        RECT  3.755 -0.250 4.015 0.755 ;
        RECT  2.995 -0.250 3.755 0.250 ;
        RECT  2.735 -0.250 2.995 0.945 ;
        RECT  1.535 -0.250 2.735 0.250 ;
        RECT  1.275 -0.250 1.535 0.405 ;
        RECT  0.385 -0.250 1.275 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.595 4.015 3.940 ;
        RECT  2.955 3.440 3.755 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  0.785 3.440 2.695 3.940 ;
        RECT  0.525 2.960 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.995 1.510 3.335 1.770 ;
        RECT  2.835 1.135 2.995 2.750 ;
        RECT  2.485 1.135 2.835 1.295 ;
        RECT  2.295 2.590 2.835 2.750 ;
        RECT  2.395 1.530 2.655 1.790 ;
        RECT  2.225 1.035 2.485 1.295 ;
        RECT  2.155 1.535 2.395 1.695 ;
        RECT  1.995 1.535 2.155 2.290 ;
        RECT  1.955 0.440 2.055 0.700 ;
        RECT  1.955 1.535 1.995 1.695 ;
        RECT  1.895 2.030 1.995 2.290 ;
        RECT  1.795 0.440 1.955 1.695 ;
        RECT  1.095 1.030 1.795 1.190 ;
        RECT  1.075 2.170 1.335 2.430 ;
        RECT  0.835 1.030 1.095 1.290 ;
        RECT  0.385 2.170 1.075 2.330 ;
        RECT  0.125 2.170 0.385 2.430 ;
    END
END AOI211X4

MACRO AOI211X2
    CLASS CORE ;
    FOREIGN AOI211X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.995 0.695 4.015 0.945 ;
        RECT  3.995 2.110 4.015 2.430 ;
        RECT  3.835 0.475 3.995 2.430 ;
        RECT  3.735 0.475 3.835 1.075 ;
        RECT  3.805 2.110 3.835 2.430 ;
        RECT  3.175 2.270 3.805 2.430 ;
        RECT  2.885 0.915 3.735 1.075 ;
        RECT  2.915 2.270 3.175 2.870 ;
        RECT  1.945 0.755 2.885 1.075 ;
        RECT  0.455 0.915 1.945 1.075 ;
        RECT  0.295 0.615 0.455 1.075 ;
        RECT  0.195 0.615 0.295 0.875 ;
        END
        ANTENNADIFFAREA     1.5119 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 1.305 3.655 1.645 ;
        RECT  2.525 1.305 3.395 1.465 ;
        RECT  2.265 1.305 2.525 1.755 ;
        RECT  2.175 1.305 2.265 1.580 ;
        RECT  1.965 1.290 2.175 1.580 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 1.675 3.175 2.045 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.845 1.255 1.255 1.580 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.645 1.445 1.745 1.705 ;
        RECT  1.485 1.445 1.645 1.920 ;
        RECT  0.625 1.760 1.485 1.920 ;
        RECT  0.465 1.255 0.625 1.920 ;
        RECT  0.365 1.255 0.465 1.580 ;
        RECT  0.125 1.290 0.365 1.580 ;
        END
        ANTENNAGATEAREA     0.4342 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.475 -0.250 4.140 0.250 ;
        RECT  3.215 -0.250 3.475 0.735 ;
        RECT  1.275 -0.250 3.215 0.250 ;
        RECT  1.015 -0.250 1.275 0.735 ;
        RECT  0.000 -0.250 1.015 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 3.440 4.140 3.940 ;
        RECT  1.695 3.285 1.955 3.940 ;
        RECT  0.895 3.440 1.695 3.940 ;
        RECT  0.635 2.440 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.735 2.615 3.995 3.215 ;
        RECT  2.355 3.055 3.735 3.215 ;
        RECT  2.195 2.100 2.355 3.215 ;
        RECT  2.095 2.100 2.195 2.770 ;
        RECT  1.405 2.100 2.095 2.260 ;
        RECT  1.145 2.100 1.405 2.700 ;
        RECT  0.385 2.100 1.145 2.260 ;
        RECT  0.125 2.100 0.385 2.700 ;
    END
END AOI211X2

MACRO AOI211X1
    CLASS CORE ;
    FOREIGN AOI211X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.165 2.520 2.175 2.810 ;
        RECT  2.005 0.645 2.165 2.810 ;
        RECT  1.990 0.645 2.005 0.945 ;
        RECT  1.990 2.335 2.005 2.810 ;
        RECT  1.820 0.645 1.990 0.905 ;
        RECT  1.965 2.450 1.990 2.810 ;
        RECT  1.905 2.450 1.965 2.710 ;
        RECT  1.095 0.745 1.820 0.905 ;
        RECT  0.835 0.745 1.095 1.035 ;
        END
        ANTENNADIFFAREA     0.6872 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.325 1.585 1.465 1.860 ;
        RECT  1.305 1.585 1.325 2.400 ;
        RECT  1.165 1.700 1.305 2.400 ;
        RECT  1.045 2.110 1.165 2.400 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.105 1.815 2.270 ;
        RECT  1.655 1.105 1.715 2.400 ;
        RECT  1.505 2.110 1.655 2.400 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.220 0.405 1.840 ;
        END
        ANTENNAGATEAREA     0.2028 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.455 0.985 1.860 ;
        RECT  0.585 1.455 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.2028 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 -0.250 2.300 0.250 ;
        RECT  1.245 -0.250 1.505 0.405 ;
        RECT  0.385 -0.250 1.245 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 3.440 2.300 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.075 2.650 1.335 2.910 ;
        RECT  0.385 2.650 1.075 2.810 ;
        RECT  0.125 2.145 0.385 2.810 ;
    END
END AOI211X1

MACRO AOI211XL
    CLASS CORE ;
    FOREIGN AOI211XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.165 2.110 2.175 2.585 ;
        RECT  2.155 0.950 2.165 2.585 ;
        RECT  2.140 0.950 2.155 2.660 ;
        RECT  2.005 0.850 2.140 2.660 ;
        RECT  1.880 0.850 2.005 1.110 ;
        RECT  1.965 2.110 2.005 2.660 ;
        RECT  1.895 2.400 1.965 2.660 ;
        RECT  1.690 0.880 1.880 1.110 ;
        RECT  1.095 0.950 1.690 1.110 ;
        RECT  0.835 0.850 1.095 1.110 ;
        END
        ANTENNADIFFAREA     0.4264 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.975 1.290 1.345 1.580 ;
        RECT  0.755 1.290 0.975 1.520 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 1.425 1.825 1.990 ;
        RECT  1.505 1.700 1.565 1.990 ;
        END
        ANTENNAGATEAREA     0.1040 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.405 1.770 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.765 1.035 2.215 ;
        RECT  0.585 1.700 0.795 2.215 ;
        END
        ANTENNAGATEAREA     0.1157 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.560 -0.250 2.300 0.250 ;
        RECT  1.300 -0.250 1.560 0.405 ;
        RECT  0.385 -0.250 1.300 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 3.440 2.300 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.075 2.400 1.335 2.660 ;
        RECT  0.385 2.400 1.075 2.560 ;
        RECT  0.125 2.400 0.385 2.660 ;
    END
END AOI211XL

MACRO AOI21X4
    CLASS CORE ;
    FOREIGN AOI21X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.895 2.335 4.935 3.000 ;
        RECT  4.835 2.255 4.895 3.195 ;
        RECT  4.635 1.790 4.835 3.195 ;
        RECT  4.475 1.790 4.635 1.990 ;
        RECT  3.875 2.995 4.635 3.195 ;
        RECT  4.465 1.290 4.475 1.990 ;
        RECT  4.265 1.075 4.465 1.990 ;
        RECT  3.815 1.075 4.265 1.275 ;
        RECT  3.615 2.595 3.875 3.195 ;
        RECT  3.555 0.675 3.815 1.275 ;
        RECT  2.450 1.005 3.555 1.205 ;
        RECT  2.355 0.880 2.450 1.205 ;
        RECT  2.095 0.605 2.355 1.205 ;
        RECT  0.385 1.005 2.095 1.205 ;
        RECT  0.125 0.605 0.385 1.205 ;
        END
        ANTENNADIFFAREA     1.7046 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.510 3.985 1.770 ;
        RECT  3.345 1.510 3.555 1.990 ;
        END
        ANTENNAGATEAREA     0.6435 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.075 1.700 3.095 1.990 ;
        RECT  3.070 1.510 3.075 1.990 ;
        RECT  2.885 1.425 3.070 1.990 ;
        RECT  2.815 1.425 2.885 1.770 ;
        RECT  1.115 1.425 2.815 1.585 ;
        RECT  0.855 1.425 1.115 1.685 ;
        END
        ANTENNAGATEAREA     0.7254 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.995 1.765 2.595 2.025 ;
        RECT  0.605 1.865 1.995 2.025 ;
        RECT  0.445 1.510 0.605 2.025 ;
        RECT  0.345 1.510 0.445 1.990 ;
        RECT  0.125 1.700 0.345 1.990 ;
        END
        ANTENNAGATEAREA     0.7254 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.355 -0.250 5.060 0.250 ;
        RECT  4.355 0.585 4.695 0.845 ;
        RECT  4.095 -0.250 4.355 0.845 ;
        RECT  3.275 -0.250 4.095 0.250 ;
        RECT  3.015 -0.250 3.275 0.755 ;
        RECT  1.340 -0.250 3.015 0.250 ;
        RECT  1.080 -0.250 1.340 0.735 ;
        RECT  0.000 -0.250 1.080 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 3.440 5.060 3.940 ;
        RECT  2.595 2.595 2.855 3.940 ;
        RECT  1.795 3.440 2.595 3.940 ;
        RECT  1.535 3.285 1.795 3.940 ;
        RECT  0.895 3.440 1.535 3.940 ;
        RECT  0.635 2.730 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.125 2.170 4.385 2.770 ;
        RECT  3.365 2.170 4.125 2.330 ;
        RECT  3.155 2.170 3.365 3.180 ;
        RECT  3.105 2.240 3.155 3.180 ;
        RECT  2.345 2.240 3.105 2.400 ;
        RECT  2.085 2.240 2.345 3.180 ;
        RECT  1.405 2.315 2.085 2.475 ;
        RECT  1.145 2.315 1.405 2.915 ;
        RECT  0.385 2.315 1.145 2.475 ;
        RECT  0.125 2.315 0.385 3.020 ;
    END
END AOI21X4

MACRO AOI21X2
    CLASS CORE ;
    FOREIGN AOI21X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.045 1.700 3.095 1.990 ;
        RECT  2.935 1.360 3.045 2.385 ;
        RECT  2.885 1.360 2.935 2.820 ;
        RECT  2.295 1.360 2.885 1.520 ;
        RECT  2.675 2.220 2.885 2.820 ;
        RECT  2.225 0.975 2.295 1.520 ;
        RECT  2.135 0.875 2.225 1.520 ;
        RECT  1.965 0.875 2.135 1.135 ;
        RECT  0.610 0.975 1.965 1.135 ;
        RECT  0.195 0.875 0.610 1.135 ;
        END
        ANTENNADIFFAREA     0.7966 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 1.700 2.635 2.040 ;
        END
        ANTENNAGATEAREA     0.3276 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.705 1.445 1.965 ;
        RECT  1.045 1.700 1.255 1.990 ;
        RECT  0.845 1.705 1.045 1.965 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 1.700 2.055 1.960 ;
        RECT  1.795 1.360 1.955 1.960 ;
        RECT  0.555 1.360 1.795 1.520 ;
        RECT  0.395 1.360 0.555 1.895 ;
        RECT  0.335 1.635 0.395 1.895 ;
        RECT  0.295 1.635 0.335 1.990 ;
        RECT  0.125 1.700 0.295 1.990 ;
        END
        ANTENNAGATEAREA     0.3692 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.765 -0.250 3.680 0.250 ;
        RECT  2.505 -0.250 2.765 1.180 ;
        RECT  1.335 -0.250 2.505 0.250 ;
        RECT  1.075 -0.250 1.335 0.795 ;
        RECT  0.000 -0.250 1.075 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 3.440 3.680 3.940 ;
        RECT  1.655 2.755 1.915 3.940 ;
        RECT  0.895 3.440 1.655 3.940 ;
        RECT  0.635 2.755 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.225 2.420 3.485 3.160 ;
        RECT  2.425 3.000 3.225 3.160 ;
        RECT  2.265 2.285 2.425 3.160 ;
        RECT  2.165 2.285 2.265 2.885 ;
        RECT  1.405 2.285 2.165 2.445 ;
        RECT  1.145 2.285 1.405 2.885 ;
        RECT  0.385 2.285 1.145 2.445 ;
        RECT  0.125 2.285 0.385 2.920 ;
    END
END AOI21X2

MACRO AOI21X1
    CLASS CORE ;
    FOREIGN AOI21X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 1.515 2.175 2.400 ;
        RECT  1.965 1.200 2.125 2.400 ;
        RECT  1.405 1.200 1.965 1.360 ;
        RECT  1.915 2.180 1.965 2.400 ;
        RECT  1.655 2.180 1.915 2.780 ;
        RECT  1.245 0.850 1.405 1.360 ;
        RECT  1.145 0.850 1.245 1.110 ;
        END
        ANTENNADIFFAREA     0.4820 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.540 1.715 1.990 ;
        RECT  1.315 1.540 1.505 1.800 ;
        END
        ANTENNAGATEAREA     0.1638 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.385 1.770 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.615 1.035 1.985 ;
        RECT  0.715 1.615 0.795 1.990 ;
        RECT  0.585 1.700 0.715 1.990 ;
        END
        ANTENNAGATEAREA     0.1846 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 -0.250 2.300 0.250 ;
        RECT  1.655 -0.250 1.915 1.015 ;
        RECT  0.585 -0.250 1.655 0.250 ;
        RECT  0.325 -0.250 0.585 1.015 ;
        RECT  0.000 -0.250 0.325 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 3.440 2.300 3.940 ;
        RECT  0.635 2.640 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.145 2.280 1.405 2.880 ;
        RECT  0.385 2.280 1.145 2.440 ;
        RECT  0.125 2.280 0.385 2.880 ;
    END
END AOI21X1

MACRO AOI21XL
    CLASS CORE ;
    FOREIGN AOI21XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 1.515 2.175 2.400 ;
        RECT  1.990 1.250 2.125 2.400 ;
        RECT  1.965 1.250 1.990 2.555 ;
        RECT  1.405 1.250 1.965 1.410 ;
        RECT  1.755 2.240 1.965 2.555 ;
        RECT  1.655 2.295 1.755 2.555 ;
        RECT  1.245 0.820 1.405 1.410 ;
        RECT  1.145 0.820 1.245 1.080 ;
        END
        ANTENNADIFFAREA     0.2806 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 1.605 1.715 1.990 ;
        RECT  1.505 1.600 1.575 1.990 ;
        RECT  1.315 1.600 1.505 1.860 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.385 1.770 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.935 1.675 1.035 1.935 ;
        RECT  0.795 1.420 0.935 1.935 ;
        RECT  0.775 1.290 0.795 1.935 ;
        RECT  0.585 1.290 0.775 1.580 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 -0.250 2.300 0.250 ;
        RECT  1.715 -0.250 1.975 1.070 ;
        RECT  0.585 -0.250 1.715 0.250 ;
        RECT  0.325 -0.250 0.585 1.070 ;
        RECT  0.000 -0.250 0.325 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 3.440 2.300 3.940 ;
        RECT  0.635 2.455 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.305 2.295 1.405 2.555 ;
        RECT  1.145 2.115 1.305 2.555 ;
        RECT  0.385 2.115 1.145 2.275 ;
        RECT  0.225 2.115 0.385 2.555 ;
        RECT  0.125 2.295 0.225 2.555 ;
    END
END AOI21XL

MACRO AND4X8
    CLASS CORE ;
    FOREIGN AND4X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 0.915 6.775 2.585 ;
        RECT  6.465 0.695 6.725 2.895 ;
        RECT  6.105 0.915 6.465 2.400 ;
        RECT  5.775 0.915 6.105 1.315 ;
        RECT  5.705 1.975 6.105 2.400 ;
        RECT  5.460 0.615 5.775 1.315 ;
        RECT  5.460 1.975 5.705 3.045 ;
        RECT  5.445 2.105 5.460 3.045 ;
        END
        ANTENNADIFFAREA     1.5844 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 1.325 4.940 1.585 ;
        RECT  4.675 1.325 4.835 2.740 ;
        RECT  1.825 2.580 4.675 2.740 ;
        RECT  1.665 1.955 1.825 2.740 ;
        RECT  1.565 1.955 1.665 2.400 ;
        RECT  1.505 2.110 1.565 2.400 ;
        END
        ANTENNAGATEAREA     0.5304 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.360 1.325 4.460 1.765 ;
        RECT  4.200 1.325 4.360 2.270 ;
        RECT  2.635 2.110 4.200 2.270 ;
        RECT  2.425 2.110 2.635 2.400 ;
        RECT  2.335 2.110 2.425 2.270 ;
        RECT  2.175 1.605 2.335 2.270 ;
        RECT  2.075 1.605 2.175 1.905 ;
        RECT  1.345 1.605 2.075 1.765 ;
        RECT  1.085 1.605 1.345 1.905 ;
        END
        ANTENNAGATEAREA     0.5304 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.720 1.645 3.980 1.925 ;
        RECT  2.850 1.765 3.720 1.925 ;
        RECT  2.690 1.265 2.850 1.925 ;
        RECT  2.590 1.265 2.690 1.585 ;
        RECT  0.865 1.265 2.590 1.425 ;
        RECT  0.795 1.265 0.865 1.905 ;
        RECT  0.705 1.265 0.795 1.990 ;
        RECT  0.585 1.515 0.705 1.990 ;
        END
        ANTENNAGATEAREA     0.5304 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.265 1.325 3.365 1.585 ;
        RECT  3.105 0.925 3.265 1.585 ;
        RECT  0.385 0.925 3.105 1.085 ;
        RECT  0.225 0.925 0.385 1.595 ;
        RECT  0.125 1.290 0.225 1.595 ;
        END
        ANTENNAGATEAREA     0.5304 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 -0.250 7.360 0.250 ;
        RECT  6.975 -0.250 7.235 1.275 ;
        RECT  6.215 -0.250 6.975 0.250 ;
        RECT  5.955 -0.250 6.215 0.735 ;
        RECT  5.140 -0.250 5.955 0.250 ;
        RECT  4.880 -0.250 5.140 0.805 ;
        RECT  1.855 -0.250 4.880 0.250 ;
        RECT  1.595 -0.250 1.855 0.405 ;
        RECT  0.000 -0.250 1.595 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 3.440 7.360 3.940 ;
        RECT  6.975 2.255 7.235 3.940 ;
        RECT  6.215 3.440 6.975 3.940 ;
        RECT  5.955 2.595 6.215 3.940 ;
        RECT  5.160 3.440 5.955 3.940 ;
        RECT  4.900 3.285 5.160 3.940 ;
        RECT  4.080 3.440 4.900 3.940 ;
        RECT  3.820 3.285 4.080 3.940 ;
        RECT  3.000 3.440 3.820 3.940 ;
        RECT  2.740 3.285 3.000 3.940 ;
        RECT  1.915 3.440 2.740 3.940 ;
        RECT  1.655 3.285 1.915 3.940 ;
        RECT  0.865 3.440 1.655 3.940 ;
        RECT  0.605 2.540 0.865 3.940 ;
        RECT  0.000 3.440 0.605 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.280 1.520 5.875 1.780 ;
        RECT  5.175 0.985 5.280 1.925 ;
        RECT  5.120 0.985 5.175 3.080 ;
        RECT  3.655 0.985 5.120 1.145 ;
        RECT  5.015 1.765 5.120 3.080 ;
        RECT  4.620 2.920 5.015 3.080 ;
        RECT  4.360 2.920 4.620 3.195 ;
        RECT  3.540 2.920 4.360 3.080 ;
        RECT  3.495 0.585 3.655 1.145 ;
        RECT  3.280 2.920 3.540 3.195 ;
        RECT  0.125 0.585 3.495 0.745 ;
        RECT  2.460 2.920 3.280 3.080 ;
        RECT  2.200 2.920 2.460 3.195 ;
        RECT  1.375 2.920 2.200 3.080 ;
        RECT  1.115 2.580 1.375 3.180 ;
    END
END AND4X8

MACRO AND4X6
    CLASS CORE ;
    FOREIGN AND4X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.815 1.515 5.855 2.585 ;
        RECT  5.535 1.290 5.815 2.895 ;
        RECT  5.515 0.695 5.535 2.895 ;
        RECT  5.370 0.695 5.515 2.400 ;
        RECT  5.255 0.695 5.370 2.285 ;
        RECT  4.835 0.885 5.255 2.285 ;
        RECT  4.710 0.885 4.835 2.915 ;
        RECT  4.495 0.885 4.710 1.185 ;
        RECT  4.535 1.975 4.710 2.915 ;
        RECT  4.190 0.495 4.495 1.185 ;
        END
        ANTENNADIFFAREA     1.5392 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.915 1.845 4.015 2.175 ;
        RECT  3.755 1.845 3.915 2.465 ;
        RECT  0.525 2.305 3.755 2.465 ;
        RECT  0.365 1.495 0.525 2.465 ;
        RECT  0.265 1.495 0.365 1.990 ;
        RECT  0.125 1.700 0.265 1.990 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.535 1.290 3.555 1.700 ;
        RECT  3.275 1.290 3.535 1.995 ;
        RECT  2.785 1.290 3.275 1.450 ;
        RECT  2.625 0.950 2.785 1.450 ;
        RECT  1.325 0.950 2.625 1.110 ;
        RECT  1.165 0.950 1.325 1.885 ;
        RECT  1.070 1.105 1.165 1.885 ;
        RECT  1.045 1.105 1.070 1.985 ;
        RECT  0.775 1.725 1.045 1.985 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.700 3.095 1.990 ;
        RECT  2.725 1.730 2.885 1.990 ;
        RECT  2.515 1.730 2.725 2.125 ;
        RECT  1.815 1.965 2.515 2.125 ;
        RECT  1.555 1.805 1.815 2.125 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 1.465 2.295 1.745 ;
        RECT  1.715 1.465 2.035 1.625 ;
        RECT  1.505 1.290 1.715 1.625 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.005 -0.250 5.980 0.250 ;
        RECT  4.745 -0.250 5.005 0.705 ;
        RECT  3.920 -0.250 4.745 0.250 ;
        RECT  3.660 -0.250 3.920 0.745 ;
        RECT  0.850 -0.250 3.660 0.250 ;
        RECT  0.590 -0.250 0.850 1.295 ;
        RECT  0.000 -0.250 0.590 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.305 3.440 5.980 3.940 ;
        RECT  5.045 2.595 5.305 3.940 ;
        RECT  4.220 3.440 5.045 3.940 ;
        RECT  3.960 3.285 4.220 3.940 ;
        RECT  3.420 3.440 3.960 3.940 ;
        RECT  3.160 3.285 3.420 3.940 ;
        RECT  2.360 3.440 3.160 3.940 ;
        RECT  2.100 2.985 2.360 3.940 ;
        RECT  1.300 3.440 2.100 3.940 ;
        RECT  1.040 3.285 1.300 3.940 ;
        RECT  0.385 3.440 1.040 3.940 ;
        RECT  0.125 2.745 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.355 1.455 4.495 1.715 ;
        RECT  4.195 1.455 4.355 2.805 ;
        RECT  3.895 1.455 4.195 1.615 ;
        RECT  3.820 2.645 4.195 2.805 ;
        RECT  3.735 0.950 3.895 1.615 ;
        RECT  3.560 2.645 3.820 2.905 ;
        RECT  3.325 0.950 3.735 1.110 ;
        RECT  2.870 2.645 3.560 2.805 ;
        RECT  3.165 0.610 3.325 1.110 ;
        RECT  2.295 0.610 3.165 0.770 ;
        RECT  2.610 2.645 2.870 2.905 ;
        RECT  1.850 2.645 2.610 2.805 ;
        RECT  2.035 0.510 2.295 0.770 ;
        RECT  1.590 2.645 1.850 2.905 ;
        RECT  0.895 2.645 1.590 2.805 ;
        RECT  0.635 2.645 0.895 2.905 ;
    END
END AND4X6

MACRO AND4X4
    CLASS CORE ;
    FOREIGN AND4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.235 1.035 4.475 2.215 ;
        RECT  3.870 1.035 4.235 1.275 ;
        RECT  3.870 1.975 4.235 2.215 ;
        RECT  3.610 0.675 3.870 1.275 ;
        RECT  3.610 1.975 3.870 2.915 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.920 1.295 3.080 2.480 ;
        RECT  2.890 1.295 2.920 1.555 ;
        RECT  2.375 2.320 2.920 2.480 ;
        RECT  2.215 2.320 2.375 2.740 ;
        RECT  0.420 2.580 2.215 2.740 ;
        RECT  0.420 1.305 0.515 1.565 ;
        RECT  0.260 1.305 0.420 2.740 ;
        RECT  0.255 1.305 0.260 2.585 ;
        RECT  0.125 1.515 0.255 2.585 ;
        END
        ANTENNAGATEAREA     0.2652 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.975 2.710 2.135 ;
        RECT  2.590 1.515 2.635 2.135 ;
        RECT  2.430 1.270 2.590 2.135 ;
        RECT  2.425 1.270 2.430 1.990 ;
        RECT  2.270 1.270 2.425 1.430 ;
        RECT  2.110 1.075 2.270 1.430 ;
        RECT  0.865 1.075 2.110 1.235 ;
        RECT  0.705 1.075 0.865 2.125 ;
        RECT  0.605 1.865 0.705 2.125 ;
        END
        ANTENNAGATEAREA     0.2652 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.880 1.880 2.140 2.140 ;
        RECT  1.715 1.980 1.880 2.140 ;
        RECT  1.555 1.980 1.715 2.400 ;
        RECT  1.505 2.110 1.555 2.400 ;
        END
        ANTENNAGATEAREA     0.2652 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.400 1.445 1.660 1.705 ;
        RECT  1.255 1.545 1.400 1.705 ;
        RECT  1.095 1.545 1.255 1.990 ;
        RECT  1.045 1.700 1.095 1.990 ;
        END
        ANTENNAGATEAREA     0.2652 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 -0.250 4.600 0.250 ;
        RECT  4.150 -0.250 4.410 0.835 ;
        RECT  3.300 -0.250 4.150 0.250 ;
        RECT  3.040 -0.250 3.300 0.750 ;
        RECT  0.390 -0.250 3.040 0.250 ;
        RECT  0.130 -0.250 0.390 0.945 ;
        RECT  0.000 -0.250 0.130 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 3.440 4.600 3.940 ;
        RECT  4.150 2.505 4.410 3.940 ;
        RECT  3.360 3.440 4.150 3.940 ;
        RECT  3.100 3.005 3.360 3.940 ;
        RECT  2.100 3.440 3.100 3.940 ;
        RECT  1.840 3.285 2.100 3.940 ;
        RECT  1.020 3.440 1.840 3.940 ;
        RECT  0.760 2.945 1.020 3.940 ;
        RECT  0.000 3.440 0.760 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.430 1.495 3.880 1.755 ;
        RECT  3.270 0.930 3.430 2.825 ;
        RECT  2.815 0.930 3.270 1.090 ;
        RECT  2.815 2.665 3.270 2.825 ;
        RECT  2.655 0.635 2.815 1.090 ;
        RECT  2.555 2.665 2.815 3.080 ;
        RECT  1.830 0.635 2.655 0.795 ;
        RECT  1.560 2.920 2.555 3.080 ;
        RECT  1.570 0.635 1.830 0.895 ;
        RECT  1.300 2.920 1.560 3.195 ;
    END
END AND4X4

MACRO AND4X2
    CLASS CORE ;
    FOREIGN AND4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 0.695 3.095 2.895 ;
        RECT  2.885 0.695 2.910 1.700 ;
        RECT  2.835 1.955 2.910 2.895 ;
        RECT  2.835 0.695 2.885 1.295 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.370 1.985 1.650 ;
        RECT  1.505 1.290 1.715 1.650 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.990 2.520 2.175 2.810 ;
        RECT  1.965 2.520 1.990 3.045 ;
        RECT  1.655 2.650 1.965 3.045 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 2.790 1.035 3.215 ;
        RECT  0.690 2.790 0.795 3.220 ;
        RECT  0.585 2.930 0.690 3.220 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.535 1.705 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 -0.250 3.220 0.250 ;
        RECT  2.295 -0.250 2.555 0.745 ;
        RECT  0.000 -0.250 2.295 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.535 3.440 3.220 3.940 ;
        RECT  2.375 2.215 2.535 3.940 ;
        RECT  2.265 3.285 2.375 3.940 ;
        RECT  1.475 3.440 2.265 3.940 ;
        RECT  1.215 2.215 1.475 3.940 ;
        RECT  0.385 3.440 1.215 3.940 ;
        RECT  0.125 2.215 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.605 1.510 2.655 1.770 ;
        RECT  2.445 0.925 2.605 2.035 ;
        RECT  0.715 0.925 2.445 1.085 ;
        RECT  2.015 1.875 2.445 2.035 ;
        RECT  1.755 1.875 2.015 2.290 ;
        RECT  0.925 1.875 1.755 2.035 ;
        RECT  0.765 1.875 0.925 2.455 ;
        RECT  0.665 2.195 0.765 2.455 ;
        RECT  0.455 0.825 0.715 1.085 ;
    END
END AND4X2

MACRO AND4X1
    CLASS CORE ;
    FOREIGN AND4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.105 2.635 2.175 ;
        RECT  2.425 0.910 2.585 2.320 ;
        RECT  2.215 0.910 2.425 1.170 ;
        RECT  2.305 2.060 2.425 2.320 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.170 2.520 2.175 2.810 ;
        RECT  1.965 2.520 2.170 2.820 ;
        RECT  1.785 2.620 1.965 2.820 ;
        RECT  1.525 2.620 1.785 2.880 ;
        END
        ANTENNAGATEAREA     0.0715 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.670 1.395 1.930 ;
        RECT  1.095 1.290 1.255 1.930 ;
        RECT  1.045 1.290 1.095 1.765 ;
        END
        ANTENNAGATEAREA     0.0715 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.335 0.800 1.990 ;
        END
        ANTENNAGATEAREA     0.0715 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.330 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0715 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 -0.250 2.760 0.250 ;
        RECT  1.675 -0.250 1.935 0.745 ;
        RECT  0.000 -0.250 1.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.225 3.440 2.760 3.940 ;
        RECT  1.965 3.000 2.225 3.940 ;
        RECT  0.920 3.440 1.965 3.940 ;
        RECT  0.320 2.880 0.920 3.940 ;
        RECT  0.000 3.440 0.320 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.750 1.350 2.185 1.610 ;
        RECT  1.590 0.950 1.750 2.340 ;
        RECT  0.425 0.950 1.590 1.110 ;
        RECT  1.585 2.180 1.590 2.340 ;
        RECT  1.325 2.180 1.585 2.440 ;
        RECT  0.570 2.180 1.325 2.340 ;
        RECT  0.310 2.180 0.570 2.440 ;
        RECT  0.165 0.820 0.425 1.110 ;
    END
END AND4X1

MACRO AND4XL
    CLASS CORE ;
    FOREIGN AND4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.105 2.635 2.175 ;
        RECT  2.425 0.745 2.585 2.320 ;
        RECT  2.245 0.745 2.425 1.005 ;
        RECT  2.305 2.060 2.425 2.320 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.170 2.520 2.175 2.810 ;
        RECT  1.965 2.520 2.170 2.820 ;
        RECT  1.785 2.620 1.965 2.820 ;
        RECT  1.525 2.620 1.785 2.880 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.690 1.395 1.950 ;
        RECT  1.095 1.290 1.255 1.950 ;
        RECT  1.045 1.290 1.095 1.765 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.335 0.800 1.895 ;
        RECT  0.585 1.335 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.330 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 -0.250 2.760 0.250 ;
        RECT  1.675 -0.250 1.935 0.745 ;
        RECT  0.000 -0.250 1.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.225 3.440 2.760 3.940 ;
        RECT  1.965 3.000 2.225 3.940 ;
        RECT  0.920 3.440 1.965 3.940 ;
        RECT  0.320 2.880 0.920 3.940 ;
        RECT  0.000 3.440 0.320 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.750 1.370 2.185 1.630 ;
        RECT  1.590 0.950 1.750 2.340 ;
        RECT  0.390 0.950 1.590 1.110 ;
        RECT  1.585 2.180 1.590 2.340 ;
        RECT  1.325 2.180 1.585 2.440 ;
        RECT  0.570 2.180 1.325 2.340 ;
        RECT  0.310 2.180 0.570 2.440 ;
        RECT  0.130 0.745 0.390 1.110 ;
    END
END AND4XL

MACRO AND3X8
    CLASS CORE ;
    FOREIGN AND3X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.800 1.515 5.855 2.585 ;
        RECT  5.540 1.265 5.800 2.925 ;
        RECT  5.185 1.265 5.540 1.990 ;
        RECT  4.925 0.695 5.185 1.990 ;
        RECT  4.780 0.975 4.925 1.990 ;
        RECT  4.520 0.975 4.780 2.920 ;
        RECT  4.105 0.975 4.520 1.990 ;
        RECT  3.910 0.630 4.105 1.990 ;
        RECT  3.845 0.630 3.910 1.230 ;
        END
        ANTENNADIFFAREA     1.6082 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.190 1.840 3.290 2.100 ;
        RECT  3.030 1.840 3.190 2.455 ;
        RECT  0.850 2.295 3.030 2.455 ;
        RECT  0.690 1.580 0.850 2.455 ;
        RECT  0.590 1.580 0.690 2.175 ;
        RECT  0.585 1.700 0.590 2.175 ;
        END
        ANTENNAGATEAREA     0.5200 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.935 2.790 2.115 ;
        RECT  2.425 1.700 2.635 2.115 ;
        RECT  1.400 1.955 2.425 2.115 ;
        RECT  1.145 1.935 1.400 2.115 ;
        RECT  1.140 1.935 1.145 2.095 ;
        END
        ANTENNAGATEAREA     0.5200 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 1.615 2.240 1.775 ;
        RECT  1.965 1.290 2.175 1.775 ;
        RECT  1.640 1.515 1.965 1.775 ;
        END
        ANTENNAGATEAREA     0.5200 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.725 -0.250 6.440 0.250 ;
        RECT  5.465 -0.250 5.725 1.085 ;
        RECT  4.645 -0.250 5.465 0.250 ;
        RECT  4.385 -0.250 4.645 0.795 ;
        RECT  3.430 -0.250 4.385 0.250 ;
        RECT  3.170 -0.250 3.430 1.135 ;
        RECT  0.825 -0.250 3.170 0.250 ;
        RECT  0.565 -0.250 0.825 1.145 ;
        RECT  0.000 -0.250 0.565 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.310 3.440 6.440 3.940 ;
        RECT  6.050 2.215 6.310 3.940 ;
        RECT  5.290 3.440 6.050 3.940 ;
        RECT  5.030 2.215 5.290 3.940 ;
        RECT  4.240 3.440 5.030 3.940 ;
        RECT  3.980 2.550 4.240 3.940 ;
        RECT  2.600 3.440 3.980 3.940 ;
        RECT  2.340 2.985 2.600 3.940 ;
        RECT  1.530 3.440 2.340 3.940 ;
        RECT  1.270 3.285 1.530 3.940 ;
        RECT  0.450 3.440 1.270 3.940 ;
        RECT  0.190 2.550 0.450 3.940 ;
        RECT  0.000 3.440 0.190 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.655 1.410 3.730 1.670 ;
        RECT  3.495 1.410 3.655 2.795 ;
        RECT  2.975 1.410 3.495 1.570 ;
        RECT  3.130 2.635 3.495 2.795 ;
        RECT  2.870 2.635 3.130 2.895 ;
        RECT  2.815 0.930 2.975 1.570 ;
        RECT  2.070 2.635 2.870 2.795 ;
        RECT  2.100 0.930 2.815 1.090 ;
        RECT  1.840 0.490 2.100 1.090 ;
        RECT  1.810 2.635 2.070 2.895 ;
        RECT  0.990 2.635 1.810 2.795 ;
        RECT  0.730 2.635 0.990 2.895 ;
    END
END AND3X8

MACRO AND3X6
    CLASS CORE ;
    FOREIGN AND3X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.675 0.695 4.935 2.915 ;
        RECT  3.955 1.265 4.675 2.035 ;
        RECT  3.680 0.695 3.955 2.945 ;
        RECT  3.550 0.695 3.680 1.330 ;
        RECT  3.595 1.945 3.680 2.945 ;
        END
        ANTENNADIFFAREA     1.5360 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.325 3.015 1.665 ;
        RECT  2.275 1.325 2.855 1.485 ;
        RECT  2.115 0.950 2.275 1.485 ;
        RECT  1.325 0.950 2.115 1.110 ;
        RECT  1.165 0.950 1.325 1.455 ;
        RECT  0.795 1.295 1.165 1.455 ;
        RECT  0.745 1.290 0.795 1.580 ;
        RECT  0.585 1.290 0.745 1.585 ;
        RECT  0.485 1.295 0.585 1.585 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.700 2.635 1.990 ;
        RECT  2.425 1.665 2.585 1.990 ;
        RECT  2.325 1.665 2.425 1.925 ;
        RECT  1.280 1.765 2.325 1.925 ;
        RECT  1.020 1.635 1.280 1.925 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.290 1.935 1.580 ;
        END
        ANTENNAGATEAREA     0.3926 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.395 -0.250 5.060 0.250 ;
        RECT  4.135 -0.250 4.395 1.085 ;
        RECT  3.265 -0.250 4.135 0.250 ;
        RECT  3.005 -0.250 3.265 0.755 ;
        RECT  0.975 -0.250 3.005 0.250 ;
        RECT  0.715 -0.250 0.975 1.075 ;
        RECT  0.000 -0.250 0.715 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.395 3.440 5.060 3.940 ;
        RECT  4.135 2.215 4.395 3.940 ;
        RECT  3.305 3.440 4.135 3.940 ;
        RECT  3.045 3.285 3.305 3.940 ;
        RECT  2.340 3.440 3.045 3.940 ;
        RECT  2.080 3.285 2.340 3.940 ;
        RECT  1.530 3.440 2.080 3.940 ;
        RECT  1.270 3.285 1.530 3.940 ;
        RECT  0.470 3.440 1.270 3.940 ;
        RECT  0.210 2.255 0.470 3.940 ;
        RECT  0.000 3.440 0.210 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.370 1.510 3.500 1.770 ;
        RECT  3.210 0.980 3.370 2.350 ;
        RECT  2.785 0.980 3.210 1.140 ;
        RECT  2.890 2.190 3.210 2.350 ;
        RECT  2.630 2.190 2.890 2.790 ;
        RECT  2.625 0.610 2.785 1.140 ;
        RECT  1.930 2.190 2.630 2.350 ;
        RECT  2.105 0.610 2.625 0.770 ;
        RECT  1.845 0.510 2.105 0.770 ;
        RECT  1.670 2.190 1.930 2.790 ;
        RECT  0.980 2.190 1.670 2.350 ;
        RECT  0.720 2.190 0.980 2.790 ;
    END
END AND3X6

MACRO AND3X4
    CLASS CORE ;
    FOREIGN AND3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.625 1.170 2.635 2.585 ;
        RECT  2.555 1.095 2.625 2.585 ;
        RECT  2.550 1.095 2.555 2.945 ;
        RECT  2.425 0.695 2.550 2.945 ;
        RECT  2.290 0.695 2.425 1.295 ;
        RECT  2.295 2.005 2.425 2.945 ;
        END
        ANTENNADIFFAREA     0.8268 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.345 1.290 1.715 1.670 ;
        END
        ANTENNAGATEAREA     0.2418 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 1.290 1.155 1.685 ;
        RECT  0.585 1.290 0.895 1.580 ;
        END
        ANTENNAGATEAREA     0.2418 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.290 0.405 1.715 ;
        END
        ANTENNAGATEAREA     0.2418 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.220 0.250 ;
        RECT  2.835 -0.250 3.095 1.155 ;
        RECT  1.985 -0.250 2.835 0.250 ;
        RECT  1.725 -0.250 1.985 0.750 ;
        RECT  0.000 -0.250 1.725 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.220 3.940 ;
        RECT  2.835 2.215 3.095 3.940 ;
        RECT  2.005 3.440 2.835 3.940 ;
        RECT  1.745 2.510 2.005 3.940 ;
        RECT  0.925 3.440 1.745 3.940 ;
        RECT  0.665 2.235 0.925 3.940 ;
        RECT  0.000 3.440 0.665 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.085 1.510 2.245 1.770 ;
        RECT  1.925 0.950 2.085 2.055 ;
        RECT  0.505 0.950 1.925 1.110 ;
        RECT  1.465 1.895 1.925 2.055 ;
        RECT  1.205 1.895 1.465 2.915 ;
        RECT  0.385 1.895 1.205 2.055 ;
        RECT  0.245 0.475 0.505 1.110 ;
        RECT  0.175 1.895 0.385 2.915 ;
        RECT  0.125 1.975 0.175 2.915 ;
    END
END AND3X4

MACRO AND3X2
    CLASS CORE ;
    FOREIGN AND3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.015 0.695 2.175 2.915 ;
        RECT  1.915 0.695 2.015 1.295 ;
        RECT  1.915 1.975 2.015 2.915 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.310 1.350 1.570 ;
        RECT  1.070 1.310 1.255 2.400 ;
        RECT  1.045 1.580 1.070 2.400 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.575 0.855 1.835 ;
        RECT  0.595 1.290 0.795 1.835 ;
        RECT  0.585 1.290 0.595 1.700 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.375 2.155 ;
        RECT  0.115 1.895 0.125 2.155 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 -0.250 2.300 0.250 ;
        RECT  1.305 -0.250 1.565 0.770 ;
        RECT  0.000 -0.250 1.305 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.580 3.440 2.300 3.940 ;
        RECT  0.640 3.285 1.580 3.940 ;
        RECT  0.000 3.440 0.640 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.690 1.535 1.830 1.795 ;
        RECT  1.530 0.950 1.690 2.885 ;
        RECT  0.385 0.950 1.530 1.110 ;
        RECT  1.265 2.725 1.530 2.885 ;
        RECT  1.005 2.725 1.265 2.985 ;
        RECT  0.385 2.725 1.005 2.885 ;
        RECT  0.125 0.850 0.385 1.110 ;
        RECT  0.225 2.725 0.385 3.195 ;
        RECT  0.125 3.035 0.225 3.195 ;
    END
END AND3X2

MACRO AND3X1
    CLASS CORE ;
    FOREIGN AND3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.970 0.705 2.175 3.160 ;
        RECT  1.960 0.705 1.970 3.260 ;
        RECT  1.855 0.705 1.960 0.965 ;
        RECT  1.370 3.000 1.960 3.260 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 1.675 1.440 1.935 ;
        RECT  1.255 1.675 1.280 1.835 ;
        RECT  1.095 1.290 1.255 1.835 ;
        RECT  1.045 1.290 1.095 1.580 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 0.435 1.065 0.715 ;
        RECT  0.585 0.435 0.795 0.760 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.620 0.585 2.030 ;
        END
        ANTENNAGATEAREA     0.0663 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 -0.250 2.300 0.250 ;
        RECT  1.315 -0.250 1.575 0.750 ;
        RECT  0.000 -0.250 1.315 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.950 3.440 2.300 3.940 ;
        RECT  0.690 2.675 0.950 3.940 ;
        RECT  0.000 3.440 0.690 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.630 1.145 1.780 2.275 ;
        RECT  1.620 0.950 1.630 2.275 ;
        RECT  1.470 0.950 1.620 1.305 ;
        RECT  1.040 2.115 1.620 2.275 ;
        RECT  0.385 0.950 1.470 1.110 ;
        RECT  0.880 2.115 1.040 2.495 ;
        RECT  0.440 2.335 0.880 2.495 ;
        RECT  0.280 2.335 0.440 2.860 ;
        RECT  0.125 0.950 0.385 1.295 ;
        RECT  0.180 2.600 0.280 2.860 ;
    END
END AND3X1

MACRO AND3XL
    CLASS CORE ;
    FOREIGN AND3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 0.910 2.185 2.745 ;
        RECT  2.025 0.910 2.175 3.060 ;
        RECT  1.965 0.910 2.025 1.355 ;
        RECT  1.965 2.520 2.025 3.060 ;
        RECT  1.915 2.800 1.965 3.060 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.605 1.290 1.715 1.580 ;
        RECT  1.505 1.290 1.605 1.860 ;
        RECT  1.395 1.355 1.505 1.860 ;
        RECT  1.345 1.600 1.395 1.860 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.495 0.810 2.145 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.400 0.380 2.105 ;
        RECT  0.120 1.400 0.125 1.765 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 -0.250 2.300 0.250 ;
        RECT  1.185 -0.250 1.445 0.770 ;
        RECT  0.000 -0.250 1.185 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.735 3.440 2.300 3.940 ;
        RECT  1.735 2.040 1.845 2.300 ;
        RECT  1.575 2.040 1.735 3.940 ;
        RECT  1.320 3.440 1.575 3.940 ;
        RECT  1.320 2.800 1.395 3.060 ;
        RECT  1.060 2.800 1.320 3.940 ;
        RECT  0.795 2.800 1.060 3.060 ;
        RECT  0.000 3.440 1.060 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.785 0.570 1.975 0.730 ;
        RECT  1.625 0.570 1.785 1.110 ;
        RECT  1.165 0.950 1.625 1.110 ;
        RECT  1.165 2.040 1.275 2.300 ;
        RECT  1.005 0.950 1.165 2.485 ;
        RECT  0.385 0.950 1.005 1.110 ;
        RECT  0.385 2.325 1.005 2.485 ;
        RECT  0.125 0.950 0.385 1.220 ;
        RECT  0.225 2.325 0.385 3.060 ;
        RECT  0.125 2.800 0.225 3.060 ;
    END
END AND3XL

MACRO AND2X8
    CLASS CORE ;
    FOREIGN AND2X8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 1.105 4.015 2.175 ;
        RECT  3.865 0.695 3.965 2.175 ;
        RECT  3.705 0.695 3.865 2.915 ;
        RECT  3.605 0.915 3.705 2.915 ;
        RECT  3.345 0.915 3.605 2.315 ;
        RECT  2.575 0.915 3.345 1.300 ;
        RECT  2.785 1.915 3.345 2.315 ;
        RECT  2.525 1.915 2.785 2.915 ;
        END
        ANTENNADIFFAREA     1.6990 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.615 1.600 1.875 1.975 ;
        RECT  0.510 1.815 1.615 1.975 ;
        RECT  0.335 1.570 0.510 1.975 ;
        RECT  0.250 1.570 0.335 1.990 ;
        RECT  0.125 1.700 0.250 1.990 ;
        END
        ANTENNAGATEAREA     0.4732 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 1.200 1.255 1.630 ;
        END
        ANTENNAGATEAREA     0.4732 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 -0.250 4.600 0.250 ;
        RECT  4.215 -0.250 4.475 1.075 ;
        RECT  3.455 -0.250 4.215 0.250 ;
        RECT  3.195 -0.250 3.455 0.735 ;
        RECT  2.195 -0.250 3.195 0.250 ;
        RECT  1.935 -0.250 2.195 1.055 ;
        RECT  0.385 -0.250 1.935 0.250 ;
        RECT  0.125 -0.250 0.385 1.075 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 3.440 4.600 3.940 ;
        RECT  4.145 2.535 4.405 3.940 ;
        RECT  3.325 3.440 4.145 3.940 ;
        RECT  3.065 2.535 3.325 3.940 ;
        RECT  2.275 3.440 3.065 3.940 ;
        RECT  2.015 2.495 2.275 3.940 ;
        RECT  1.985 3.285 2.015 3.940 ;
        RECT  1.185 3.440 1.985 3.940 ;
        RECT  0.925 3.285 1.185 3.940 ;
        RECT  0.385 3.440 0.925 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.275 1.520 3.165 1.680 ;
        RECT  2.115 1.260 2.275 2.315 ;
        RECT  1.595 1.260 2.115 1.420 ;
        RECT  1.735 2.155 2.115 2.315 ;
        RECT  1.475 2.155 1.735 2.755 ;
        RECT  1.435 0.860 1.595 1.420 ;
        RECT  0.785 2.155 1.475 2.315 ;
        RECT  1.205 0.860 1.435 1.020 ;
        RECT  0.945 0.760 1.205 1.020 ;
        RECT  0.525 2.155 0.785 2.755 ;
    END
END AND2X8

MACRO AND2X6
    CLASS CORE ;
    FOREIGN AND2X6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.865 1.290 4.015 2.585 ;
        RECT  3.815 1.030 3.865 2.970 ;
        RECT  3.605 0.695 3.815 2.970 ;
        RECT  3.555 0.695 3.605 2.400 ;
        RECT  3.530 1.030 3.555 2.400 ;
        RECT  2.910 1.030 3.530 2.335 ;
        RECT  2.885 1.030 2.910 2.400 ;
        RECT  2.735 1.030 2.885 1.335 ;
        RECT  2.785 2.030 2.885 2.400 ;
        RECT  2.525 2.030 2.785 2.970 ;
        RECT  2.475 0.695 2.735 1.335 ;
        END
        ANTENNADIFFAREA     1.5264 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.665 1.625 1.925 1.955 ;
        RECT  0.510 1.795 1.665 1.955 ;
        RECT  0.335 1.535 0.510 1.955 ;
        RECT  0.250 1.535 0.335 1.990 ;
        RECT  0.125 1.700 0.250 1.990 ;
        END
        ANTENNAGATEAREA     0.3640 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.360 1.375 1.615 ;
        RECT  1.045 1.290 1.255 1.615 ;
        RECT  0.775 1.360 1.045 1.615 ;
        END
        ANTENNAGATEAREA     0.3640 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.275 -0.250 4.140 0.250 ;
        RECT  3.015 -0.250 3.275 0.805 ;
        RECT  2.195 -0.250 3.015 0.250 ;
        RECT  1.935 -0.250 2.195 0.975 ;
        RECT  0.385 -0.250 1.935 0.250 ;
        RECT  0.125 -0.250 0.385 1.275 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.325 3.440 4.140 3.940 ;
        RECT  3.065 2.610 3.325 3.940 ;
        RECT  2.275 3.440 3.065 3.940 ;
        RECT  1.985 2.610 2.275 3.940 ;
        RECT  1.185 3.440 1.985 3.940 ;
        RECT  0.925 3.285 1.185 3.940 ;
        RECT  0.385 3.440 0.925 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.275 1.555 2.565 1.815 ;
        RECT  2.115 1.265 2.275 2.295 ;
        RECT  1.715 1.265 2.115 1.425 ;
        RECT  1.735 2.135 2.115 2.295 ;
        RECT  1.475 2.135 1.735 2.735 ;
        RECT  1.555 0.935 1.715 1.425 ;
        RECT  1.275 0.935 1.555 1.095 ;
        RECT  0.785 2.135 1.475 2.295 ;
        RECT  1.015 0.835 1.275 1.095 ;
        RECT  0.525 2.135 0.785 2.735 ;
    END
END AND2X6

MACRO AND2X4
    CLASS CORE ;
    FOREIGN AND2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 1.700 2.175 2.400 ;
        RECT  1.955 1.700 1.975 2.895 ;
        RECT  1.785 0.850 1.955 2.895 ;
        RECT  1.715 0.495 1.785 2.895 ;
        RECT  1.525 0.495 1.715 1.095 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.655 1.065 1.990 ;
        END
        ANTENNAGATEAREA     0.2366 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.520 0.385 2.040 ;
        END
        ANTENNAGATEAREA     0.2366 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.415 -0.250 2.760 0.250 ;
        RECT  2.155 -0.250 2.415 1.135 ;
        RECT  1.235 -0.250 2.155 0.250 ;
        RECT  0.975 -0.250 1.235 1.095 ;
        RECT  0.000 -0.250 0.975 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.515 3.440 2.760 3.940 ;
        RECT  2.255 2.580 2.515 3.940 ;
        RECT  1.435 3.440 2.255 3.940 ;
        RECT  1.175 2.555 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.290 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.450 1.565 1.500 1.825 ;
        RECT  1.290 1.275 1.450 2.370 ;
        RECT  0.725 1.275 1.290 1.435 ;
        RECT  0.895 2.210 1.290 2.370 ;
        RECT  0.635 2.210 0.895 2.890 ;
        RECT  0.565 1.100 0.725 1.435 ;
        RECT  0.385 1.100 0.565 1.260 ;
        RECT  0.125 0.660 0.385 1.260 ;
    END
END AND2X4

MACRO AND2X2
    CLASS CORE ;
    FOREIGN AND2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 0.620 1.715 2.970 ;
        RECT  1.455 0.620 1.555 1.220 ;
        RECT  1.530 1.925 1.555 2.970 ;
        RECT  1.455 2.030 1.530 2.970 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.735 1.585 0.895 2.400 ;
        RECT  0.585 1.925 0.735 2.400 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.285 0.445 1.545 ;
        RECT  0.185 1.285 0.360 1.880 ;
        RECT  0.125 1.290 0.185 1.880 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.175 -0.250 1.840 0.250 ;
        RECT  0.915 -0.250 1.175 0.405 ;
        RECT  0.000 -0.250 0.915 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 1.840 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.260 1.405 1.375 1.665 ;
        RECT  1.100 1.245 1.260 2.885 ;
        RECT  0.995 1.245 1.100 1.405 ;
        RECT  0.775 2.725 1.100 2.885 ;
        RECT  0.835 0.945 0.995 1.405 ;
        RECT  0.410 0.945 0.835 1.105 ;
        RECT  0.515 2.680 0.775 2.940 ;
        RECT  0.150 0.845 0.410 1.105 ;
    END
END AND2X2

MACRO AND2X1
    CLASS CORE ;
    FOREIGN AND2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.625 0.955 1.715 2.585 ;
        RECT  1.505 0.955 1.625 2.900 ;
        RECT  1.455 0.955 1.505 1.215 ;
        RECT  1.365 2.300 1.505 2.900 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.885 0.845 2.145 ;
        RECT  0.585 1.290 0.795 2.145 ;
        END
        ANTENNAGATEAREA     0.0598 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.400 0.405 1.990 ;
        END
        ANTENNAGATEAREA     0.0598 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 -0.250 1.840 0.250 ;
        RECT  0.935 -0.250 1.195 0.405 ;
        RECT  0.000 -0.250 0.935 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.000 3.440 1.840 3.940 ;
        RECT  0.320 3.285 1.000 3.940 ;
        RECT  0.000 3.440 0.320 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.185 1.710 1.325 1.970 ;
        RECT  1.025 0.950 1.185 2.485 ;
        RECT  0.385 0.950 1.025 1.110 ;
        RECT  0.575 2.325 1.025 2.485 ;
        RECT  0.315 2.325 0.575 2.585 ;
        RECT  0.225 0.535 0.385 1.110 ;
        RECT  0.125 0.535 0.225 0.795 ;
    END
END AND2X1

MACRO AND2XL
    CLASS CORE ;
    FOREIGN AND2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.685 1.035 1.715 2.400 ;
        RECT  1.505 1.035 1.685 2.585 ;
        RECT  1.455 1.035 1.505 1.295 ;
        RECT  1.425 2.325 1.505 2.585 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.700 0.795 2.145 ;
        RECT  0.360 1.885 0.585 2.145 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.200 0.405 1.665 ;
        END
        ANTENNAGATEAREA     0.0520 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 -0.250 1.840 0.250 ;
        RECT  0.885 -0.250 1.145 0.405 ;
        RECT  0.000 -0.250 0.885 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 3.440 1.840 3.940 ;
        RECT  0.885 2.860 1.145 3.940 ;
        RECT  0.520 3.440 0.885 3.940 ;
        RECT  0.260 3.285 0.520 3.940 ;
        RECT  0.000 3.440 0.260 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.135 1.710 1.325 1.970 ;
        RECT  0.975 0.695 1.135 2.485 ;
        RECT  0.385 0.695 0.975 0.855 ;
        RECT  0.575 2.325 0.975 2.485 ;
        RECT  0.315 2.325 0.575 2.585 ;
        RECT  0.125 0.595 0.385 0.855 ;
    END
END AND2XL

MACRO HOLDX1
    CLASS CORE ;
    FOREIGN HOLDX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION INOUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 1.035 1.715 2.005 ;
        RECT  1.395 1.845 1.445 2.005 ;
        RECT  1.135 1.845 1.395 2.375 ;
        RECT  1.045 1.845 1.135 2.175 ;
        RECT  0.725 1.845 1.045 2.005 ;
        RECT  0.565 1.675 0.725 2.005 ;
        RECT  0.455 1.675 0.565 1.935 ;
        END
        ANTENNAGATEAREA     0.0494 ;
        ANTENNADIFFAREA     0.2010 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.965 -0.250 1.840 0.250 ;
        RECT  0.705 -0.250 0.965 0.745 ;
        RECT  0.000 -0.250 0.705 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.815 3.440 1.840 3.940 ;
        RECT  0.555 2.785 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.095 1.405 1.195 1.665 ;
        RECT  0.935 1.135 1.095 1.665 ;
        RECT  0.385 1.135 0.935 1.295 ;
        RECT  0.275 1.035 0.385 1.295 ;
        RECT  0.275 2.115 0.385 2.375 ;
        RECT  0.115 1.035 0.275 2.375 ;
    END
END HOLDX1

MACRO TBUFX20
    CLASS CORE ;
    FOREIGN TBUFX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  9.530 1.105 9.535 2.585 ;
        RECT  9.525 1.105 9.530 2.695 ;
        RECT  9.500 1.105 9.525 2.895 ;
        RECT  9.265 0.695 9.500 2.895 ;
        RECT  9.240 0.695 9.265 2.695 ;
        RECT  8.505 0.915 9.240 2.695 ;
        RECT  8.480 0.915 8.505 3.085 ;
        RECT  8.405 0.695 8.480 3.085 ;
        RECT  8.220 0.695 8.405 1.515 ;
        RECT  8.245 2.095 8.405 3.085 ;
        RECT  7.485 2.095 8.245 2.695 ;
        RECT  7.460 0.915 8.220 1.515 ;
        RECT  7.225 2.095 7.485 3.085 ;
        RECT  7.200 0.695 7.460 1.515 ;
        RECT  6.465 2.095 7.225 2.695 ;
        RECT  6.440 0.915 7.200 1.515 ;
        RECT  6.205 2.095 6.465 3.085 ;
        RECT  6.180 0.695 6.440 1.515 ;
        RECT  5.445 2.095 6.205 2.730 ;
        RECT  5.415 0.915 6.180 1.515 ;
        RECT  5.375 2.095 5.445 3.120 ;
        RECT  5.255 0.750 5.415 1.515 ;
        RECT  5.185 2.180 5.375 3.120 ;
        RECT  5.155 0.750 5.255 1.010 ;
        END
        ANTENNADIFFAREA     3.9404 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.110 1.355 0.370 1.990 ;
        END
        ANTENNAGATEAREA     0.5603 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.570 4.565 1.830 ;
        RECT  3.805 1.570 4.015 1.990 ;
        RECT  3.625 1.570 3.805 1.830 ;
        END
        ANTENNAGATEAREA     0.9607 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.990 -0.250 9.660 0.250 ;
        RECT  8.730 -0.250 8.990 0.735 ;
        RECT  7.970 -0.250 8.730 0.250 ;
        RECT  7.710 -0.250 7.970 0.735 ;
        RECT  6.950 -0.250 7.710 0.250 ;
        RECT  6.690 -0.250 6.950 0.735 ;
        RECT  5.925 -0.250 6.690 0.250 ;
        RECT  5.665 -0.250 5.925 0.735 ;
        RECT  4.905 -0.250 5.665 0.250 ;
        RECT  4.645 -0.250 4.905 0.735 ;
        RECT  3.885 -0.250 4.645 0.250 ;
        RECT  3.625 -0.250 3.885 1.025 ;
        RECT  1.845 -0.250 3.625 0.250 ;
        RECT  1.585 -0.250 1.845 0.930 ;
        RECT  0.850 -0.250 1.585 0.250 ;
        RECT  0.590 -0.250 0.850 0.405 ;
        RECT  0.000 -0.250 0.590 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.015 3.440 9.660 3.940 ;
        RECT  8.755 2.955 9.015 3.940 ;
        RECT  7.995 3.440 8.755 3.940 ;
        RECT  7.735 2.955 7.995 3.940 ;
        RECT  6.975 3.440 7.735 3.940 ;
        RECT  6.715 2.955 6.975 3.940 ;
        RECT  5.955 3.440 6.715 3.940 ;
        RECT  5.695 2.955 5.955 3.940 ;
        RECT  4.935 3.440 5.695 3.940 ;
        RECT  4.675 2.615 4.935 3.940 ;
        RECT  3.915 3.440 4.675 3.940 ;
        RECT  3.655 2.615 3.915 3.940 ;
        RECT  1.845 3.440 3.655 3.940 ;
        RECT  1.585 2.890 1.845 3.940 ;
        RECT  0.850 3.440 1.585 3.940 ;
        RECT  0.590 3.285 0.850 3.940 ;
        RECT  0.000 3.440 0.590 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.940 1.725 5.195 1.985 ;
        RECT  4.945 1.245 5.075 1.505 ;
        RECT  4.785 0.915 4.945 1.505 ;
        RECT  4.935 1.725 4.940 2.330 ;
        RECT  4.780 1.825 4.935 2.330 ;
        RECT  4.395 0.915 4.785 1.075 ;
        RECT  4.425 2.170 4.780 2.330 ;
        RECT  4.165 2.170 4.425 3.215 ;
        RECT  4.295 0.475 4.395 1.075 ;
        RECT  4.135 0.475 4.295 1.385 ;
        RECT  3.405 2.170 4.165 2.330 ;
        RECT  3.375 1.225 4.135 1.385 ;
        RECT  3.305 2.065 3.405 3.005 ;
        RECT  3.115 0.640 3.375 1.385 ;
        RECT  3.145 1.720 3.305 3.005 ;
        RECT  2.865 1.720 3.145 1.880 ;
        RECT  2.355 2.845 3.145 3.005 ;
        RECT  2.370 0.640 3.115 0.800 ;
        RECT  2.635 2.065 2.895 2.665 ;
        RECT  2.705 0.985 2.865 1.880 ;
        RECT  2.605 0.985 2.705 1.280 ;
        RECT  2.370 2.065 2.635 2.225 ;
        RECT  2.210 0.640 2.370 2.225 ;
        RECT  2.255 2.710 2.355 3.005 ;
        RECT  2.095 2.550 2.255 3.005 ;
        RECT  2.095 0.640 2.210 1.270 ;
        RECT  1.405 1.110 2.095 1.270 ;
        RECT  1.335 2.550 2.095 2.710 ;
        RECT  1.885 2.020 2.030 2.280 ;
        RECT  1.725 1.500 1.885 2.280 ;
        RECT  1.040 1.500 1.725 1.660 ;
        RECT  1.245 0.820 1.405 1.270 ;
        RECT  1.075 2.440 1.335 2.710 ;
        RECT  1.075 0.820 1.245 1.080 ;
        RECT  0.710 1.400 1.040 1.660 ;
        RECT  0.550 0.920 0.710 2.430 ;
        RECT  0.385 0.920 0.550 1.080 ;
        RECT  0.385 2.270 0.550 2.430 ;
        RECT  0.125 0.820 0.385 1.080 ;
        RECT  0.125 2.270 0.385 2.870 ;
    END
END TBUFX20

MACRO TBUFX16
    CLASS CORE ;
    FOREIGN TBUFX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  7.435 0.695 7.695 2.895 ;
        RECT  6.750 0.865 7.435 2.555 ;
        RECT  6.675 0.865 6.750 2.585 ;
        RECT  6.565 0.695 6.675 2.895 ;
        RECT  6.415 0.695 6.565 1.465 ;
        RECT  6.415 1.955 6.565 2.895 ;
        RECT  5.655 0.865 6.415 1.465 ;
        RECT  5.655 1.955 6.415 2.555 ;
        RECT  5.395 0.695 5.655 1.465 ;
        RECT  5.055 1.955 5.655 2.895 ;
        RECT  4.510 0.865 5.395 1.465 ;
        RECT  4.325 2.295 5.055 2.895 ;
        RECT  4.280 0.475 4.510 1.465 ;
        RECT  4.135 0.475 4.280 1.070 ;
        END
        ANTENNADIFFAREA     3.0986 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.830 0.370 2.090 ;
        RECT  0.125 1.290 0.335 2.090 ;
        RECT  0.110 1.830 0.125 2.090 ;
        END
        ANTENNAGATEAREA     0.4602 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 1.475 3.445 1.735 ;
        RECT  2.885 1.475 3.095 1.990 ;
        RECT  2.505 1.475 2.885 1.735 ;
        END
        ANTENNAGATEAREA     0.8203 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 -0.250 7.820 0.250 ;
        RECT  6.925 -0.250 7.185 0.685 ;
        RECT  6.165 -0.250 6.925 0.250 ;
        RECT  5.905 -0.250 6.165 0.685 ;
        RECT  5.060 -0.250 5.905 0.250 ;
        RECT  4.800 -0.250 5.060 0.685 ;
        RECT  3.955 -0.250 4.800 0.250 ;
        RECT  3.695 -0.250 3.955 0.735 ;
        RECT  2.935 -0.250 3.695 0.250 ;
        RECT  2.675 -0.250 2.935 0.735 ;
        RECT  0.895 -0.250 2.675 0.250 ;
        RECT  0.635 -0.250 0.895 0.770 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 3.440 7.820 3.940 ;
        RECT  6.925 2.955 7.185 3.940 ;
        RECT  6.165 3.440 6.925 3.940 ;
        RECT  5.905 2.955 6.165 3.940 ;
        RECT  4.985 3.440 5.905 3.940 ;
        RECT  4.725 3.285 4.985 3.940 ;
        RECT  4.070 3.440 4.725 3.940 ;
        RECT  3.810 2.275 4.070 3.940 ;
        RECT  3.050 3.440 3.810 3.940 ;
        RECT  2.790 2.615 3.050 3.940 ;
        RECT  0.940 3.440 2.790 3.940 ;
        RECT  0.680 3.285 0.940 3.940 ;
        RECT  0.000 3.440 0.680 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.315 1.665 4.575 2.075 ;
        RECT  3.560 1.915 4.315 2.075 ;
        RECT  3.955 1.295 4.095 1.555 ;
        RECT  3.795 1.125 3.955 1.555 ;
        RECT  3.445 1.125 3.795 1.285 ;
        RECT  3.400 1.915 3.560 3.115 ;
        RECT  3.185 0.585 3.445 1.285 ;
        RECT  3.300 2.170 3.400 3.115 ;
        RECT  2.530 2.170 3.300 2.330 ;
        RECT  2.425 1.125 3.185 1.285 ;
        RECT  2.420 2.170 2.530 2.880 ;
        RECT  2.165 0.570 2.425 1.285 ;
        RECT  2.260 1.925 2.420 2.880 ;
        RECT  2.015 3.060 2.275 3.260 ;
        RECT  1.815 1.925 2.260 2.085 ;
        RECT  1.625 2.720 2.260 2.880 ;
        RECT  1.470 0.570 2.165 0.730 ;
        RECT  1.285 3.060 2.015 3.220 ;
        RECT  1.805 2.265 1.965 2.530 ;
        RECT  1.815 1.025 1.915 1.285 ;
        RECT  1.655 1.025 1.815 2.085 ;
        RECT  1.470 2.265 1.805 2.425 ;
        RECT  1.465 2.605 1.625 2.880 ;
        RECT  1.310 0.570 1.470 2.425 ;
        RECT  1.245 2.605 1.465 2.765 ;
        RECT  1.145 0.675 1.310 1.275 ;
        RECT  1.125 2.945 1.285 3.220 ;
        RECT  0.935 2.945 1.125 3.105 ;
        RECT  0.935 1.395 0.965 1.655 ;
        RECT  0.775 1.395 0.935 3.105 ;
        RECT  0.675 1.395 0.775 1.555 ;
        RECT  0.385 2.610 0.775 2.870 ;
        RECT  0.515 0.950 0.675 1.555 ;
        RECT  0.385 0.950 0.515 1.110 ;
        RECT  0.210 0.690 0.385 1.110 ;
        RECT  0.125 2.270 0.385 2.870 ;
        RECT  0.125 0.690 0.210 0.950 ;
    END
END TBUFX16

MACRO TBUFX12
    CLASS CORE ;
    FOREIGN TBUFX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  6.260 0.695 6.315 1.355 ;
        RECT  6.265 2.335 6.315 2.585 ;
        RECT  6.005 2.125 6.265 3.065 ;
        RECT  6.000 0.520 6.260 1.505 ;
        RECT  5.855 2.125 6.005 2.805 ;
        RECT  5.855 0.880 6.000 1.505 ;
        RECT  5.830 0.880 5.855 2.805 ;
        RECT  5.245 0.905 5.830 2.805 ;
        RECT  5.240 0.905 5.245 3.065 ;
        RECT  5.185 0.520 5.240 3.065 ;
        RECT  4.980 0.520 5.185 1.505 ;
        RECT  4.985 2.125 5.185 3.065 ;
        RECT  4.820 2.125 4.985 2.895 ;
        RECT  4.910 0.880 4.980 1.505 ;
        RECT  4.290 0.905 4.910 1.505 ;
        RECT  4.035 2.295 4.820 2.895 ;
        RECT  4.170 0.495 4.290 1.505 ;
        RECT  3.935 0.495 4.170 1.135 ;
        END
        ANTENNADIFFAREA     2.3098 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 2.000 0.375 2.260 ;
        RECT  0.125 1.290 0.335 2.260 ;
        RECT  0.115 1.925 0.125 2.260 ;
        END
        ANTENNAGATEAREA     0.3419 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 1.475 3.415 1.735 ;
        RECT  2.885 1.475 3.095 1.990 ;
        RECT  2.475 1.475 2.885 1.735 ;
        END
        ANTENNAGATEAREA     0.6370 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.770 -0.250 6.900 0.250 ;
        RECT  6.510 -0.250 6.770 1.075 ;
        RECT  5.750 -0.250 6.510 0.250 ;
        RECT  5.490 -0.250 5.750 0.685 ;
        RECT  4.730 -0.250 5.490 0.250 ;
        RECT  4.470 -0.250 4.730 0.685 ;
        RECT  3.680 -0.250 4.470 0.250 ;
        RECT  3.420 -0.250 3.680 0.405 ;
        RECT  2.870 -0.250 3.420 0.250 ;
        RECT  2.610 -0.250 2.870 0.405 ;
        RECT  0.900 -0.250 2.610 0.250 ;
        RECT  0.640 -0.250 0.900 0.405 ;
        RECT  0.000 -0.250 0.640 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.255 6.775 3.940 ;
        RECT  5.755 3.440 6.515 3.940 ;
        RECT  5.495 2.985 5.755 3.940 ;
        RECT  4.695 3.440 5.495 3.940 ;
        RECT  4.435 3.285 4.695 3.940 ;
        RECT  3.745 3.440 4.435 3.940 ;
        RECT  3.485 3.285 3.745 3.940 ;
        RECT  2.795 3.440 3.485 3.940 ;
        RECT  2.535 3.285 2.795 3.940 ;
        RECT  0.820 3.440 2.535 3.940 ;
        RECT  0.560 3.285 0.820 3.940 ;
        RECT  0.000 3.440 0.560 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.215 1.685 4.520 2.075 ;
        RECT  3.435 1.915 4.215 2.075 ;
        RECT  3.755 1.315 3.990 1.575 ;
        RECT  3.595 1.135 3.755 1.575 ;
        RECT  3.270 1.135 3.595 1.295 ;
        RECT  3.275 1.915 3.435 2.915 ;
        RECT  3.085 2.260 3.275 2.915 ;
        RECT  3.010 0.925 3.270 1.295 ;
        RECT  2.395 2.260 3.085 2.420 ;
        RECT  2.290 1.135 3.010 1.295 ;
        RECT  2.285 2.215 2.395 2.815 ;
        RECT  2.130 0.430 2.290 1.295 ;
        RECT  2.135 1.475 2.285 2.815 ;
        RECT  2.125 1.475 2.135 2.765 ;
        RECT  2.030 0.430 2.130 0.730 ;
        RECT  1.880 1.475 2.125 1.635 ;
        RECT  1.115 2.605 2.125 2.765 ;
        RECT  1.480 0.570 2.030 0.730 ;
        RECT  1.380 2.265 1.885 2.425 ;
        RECT  1.720 1.090 1.880 1.635 ;
        RECT  1.620 1.090 1.720 1.350 ;
        RECT  1.375 2.945 1.635 3.235 ;
        RECT  1.380 0.430 1.480 0.730 ;
        RECT  1.220 0.430 1.380 2.425 ;
        RECT  0.715 2.945 1.375 3.105 ;
        RECT  0.715 1.530 0.890 1.790 ;
        RECT  0.555 0.920 0.715 3.105 ;
        RECT  0.385 0.920 0.555 1.080 ;
        RECT  0.165 2.610 0.555 2.870 ;
        RECT  0.125 0.820 0.385 1.080 ;
    END
END TBUFX12

MACRO TBUFX8
    CLASS CORE ;
    FOREIGN TBUFX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 0.695 4.935 2.585 ;
        RECT  4.625 0.585 4.885 3.000 ;
        RECT  3.865 1.290 4.625 1.990 ;
        RECT  3.605 0.575 3.865 3.150 ;
        END
        ANTENNADIFFAREA     1.5722 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.530 0.535 1.990 ;
        END
        ANTENNAGATEAREA     0.2301 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.255 1.545 2.605 1.705 ;
        RECT  2.095 1.545 2.255 2.735 ;
        RECT  1.965 1.700 2.095 1.990 ;
        RECT  1.325 2.575 2.095 2.735 ;
        RECT  1.165 2.035 1.325 2.735 ;
        RECT  1.065 2.035 1.165 2.295 ;
        END
        ANTENNAGATEAREA     0.4212 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 -0.250 5.520 0.250 ;
        RECT  5.135 -0.250 5.395 1.075 ;
        RECT  4.375 -0.250 5.135 0.250 ;
        RECT  4.115 -0.250 4.375 1.075 ;
        RECT  3.315 -0.250 4.115 0.250 ;
        RECT  3.055 -0.250 3.315 0.685 ;
        RECT  2.235 -0.250 3.055 0.250 ;
        RECT  1.975 -0.250 2.235 0.405 ;
        RECT  0.250 -0.250 1.975 0.250 ;
        RECT  0.355 1.030 0.615 1.290 ;
        RECT  0.250 1.030 0.355 1.190 ;
        RECT  0.090 -0.250 0.250 1.190 ;
        RECT  0.000 -0.250 0.090 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.395 3.440 5.520 3.940 ;
        RECT  5.135 2.275 5.395 3.940 ;
        RECT  4.375 3.440 5.135 3.940 ;
        RECT  4.115 2.275 4.375 3.940 ;
        RECT  3.265 3.440 4.115 3.940 ;
        RECT  3.005 2.275 3.265 3.940 ;
        RECT  0.955 3.440 3.005 3.940 ;
        RECT  0.695 3.285 0.955 3.940 ;
        RECT  0.000 3.440 0.695 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.215 0.865 3.375 1.545 ;
        RECT  2.950 1.765 3.360 2.045 ;
        RECT  2.775 0.865 3.215 1.025 ;
        RECT  2.790 1.205 2.950 2.045 ;
        RECT  1.865 1.205 2.790 1.365 ;
        RECT  2.695 1.885 2.790 2.045 ;
        RECT  2.515 0.615 2.775 1.025 ;
        RECT  2.535 1.885 2.695 3.125 ;
        RECT  2.435 2.185 2.535 3.125 ;
        RECT  1.395 0.615 2.515 0.775 ;
        RECT  1.495 2.915 2.435 3.075 ;
        RECT  1.725 2.235 1.915 2.395 ;
        RECT  1.700 0.960 1.865 1.365 ;
        RECT  1.565 1.655 1.725 2.395 ;
        RECT  1.605 0.960 1.700 1.220 ;
        RECT  1.395 1.655 1.565 1.815 ;
        RECT  1.235 2.915 1.495 3.175 ;
        RECT  1.235 0.615 1.395 1.815 ;
        RECT  1.145 1.035 1.235 1.295 ;
        RECT  0.385 2.915 1.235 3.075 ;
        RECT  0.965 1.550 1.055 1.810 ;
        RECT  0.885 0.545 0.965 1.810 ;
        RECT  0.805 0.545 0.885 2.335 ;
        RECT  0.690 0.545 0.805 0.705 ;
        RECT  0.725 1.650 0.805 2.335 ;
        RECT  0.125 2.175 0.725 2.335 ;
        RECT  0.430 0.445 0.690 0.705 ;
        RECT  0.125 2.915 0.385 3.175 ;
    END
END TBUFX8

MACRO TBUFX6
    CLASS CORE ;
    FOREIGN TBUFX6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  4.215 0.675 4.475 2.915 ;
        RECT  3.525 1.255 4.215 2.095 ;
        RECT  3.265 0.495 3.525 3.150 ;
        RECT  3.195 0.495 3.265 1.095 ;
        RECT  3.195 2.210 3.265 3.150 ;
        END
        ANTENNADIFFAREA     1.4874 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.845 0.505 2.105 ;
        RECT  0.125 1.700 0.335 2.105 ;
        END
        ANTENNAGATEAREA     0.1781 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 1.555 2.205 2.735 ;
        RECT  1.965 1.555 2.045 1.990 ;
        RECT  1.335 2.575 2.045 2.735 ;
        RECT  1.725 1.555 1.965 1.715 ;
        RECT  1.075 2.385 1.335 2.735 ;
        END
        ANTENNAGATEAREA     0.3042 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 -0.250 4.600 0.250 ;
        RECT  3.705 -0.250 3.965 1.075 ;
        RECT  2.850 -0.250 3.705 0.250 ;
        RECT  2.590 -0.250 2.850 0.405 ;
        RECT  0.265 -0.250 2.590 0.250 ;
        RECT  0.445 1.030 0.605 1.295 ;
        RECT  0.265 1.030 0.445 1.190 ;
        RECT  0.105 -0.250 0.265 1.190 ;
        RECT  0.000 -0.250 0.105 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 3.440 4.600 3.940 ;
        RECT  3.705 2.275 3.965 3.940 ;
        RECT  2.895 3.440 3.705 3.940 ;
        RECT  2.735 2.275 2.895 3.940 ;
        RECT  0.955 3.440 2.735 3.940 ;
        RECT  0.695 3.285 0.955 3.940 ;
        RECT  0.000 3.440 0.695 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.825 1.765 3.085 2.025 ;
        RECT  2.965 1.285 3.065 1.545 ;
        RECT  2.805 0.695 2.965 1.545 ;
        RECT  2.555 1.770 2.825 2.025 ;
        RECT  2.380 0.695 2.805 0.855 ;
        RECT  2.395 1.085 2.555 3.075 ;
        RECT  1.845 1.085 2.395 1.245 ;
        RECT  0.385 2.915 2.395 3.075 ;
        RECT  2.220 0.475 2.380 0.855 ;
        RECT  1.985 0.475 2.220 0.735 ;
        RECT  1.395 0.575 1.985 0.735 ;
        RECT  1.765 2.235 1.865 2.395 ;
        RECT  1.585 0.985 1.845 1.245 ;
        RECT  1.605 1.905 1.765 2.395 ;
        RECT  1.395 1.905 1.605 2.065 ;
        RECT  1.235 0.575 1.395 2.065 ;
        RECT  1.125 1.035 1.235 1.295 ;
        RECT  0.945 1.605 1.055 1.865 ;
        RECT  0.845 0.560 0.945 1.865 ;
        RECT  0.785 0.560 0.845 2.445 ;
        RECT  0.605 0.560 0.785 0.720 ;
        RECT  0.685 1.700 0.785 2.445 ;
        RECT  0.125 2.285 0.685 2.445 ;
        RECT  0.445 0.460 0.605 0.720 ;
        RECT  0.125 2.915 0.385 3.175 ;
    END
END TBUFX6

MACRO TBUFX4
    CLASS CORE ;
    FOREIGN TBUFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.290 4.015 1.990 ;
        RECT  3.555 1.510 3.805 1.770 ;
        RECT  3.505 0.695 3.555 2.585 ;
        RECT  3.245 0.575 3.505 3.030 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.600 0.505 1.860 ;
        RECT  0.125 1.600 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1326 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.945 2.260 2.400 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 -0.250 4.140 0.250 ;
        RECT  3.755 -0.250 4.015 1.075 ;
        RECT  2.795 -0.250 3.755 0.250 ;
        RECT  2.535 -0.250 2.795 1.075 ;
        RECT  0.385 -0.250 2.535 0.250 ;
        RECT  0.125 -0.250 0.385 0.855 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.275 4.015 3.940 ;
        RECT  2.795 3.440 3.755 3.940 ;
        RECT  2.535 2.275 2.795 3.940 ;
        RECT  0.385 3.440 2.535 3.940 ;
        RECT  0.125 2.920 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.995 1.265 2.735 1.425 ;
        RECT  2.730 1.775 2.735 2.035 ;
        RECT  2.475 1.605 2.730 2.035 ;
        RECT  1.775 1.605 2.475 1.765 ;
        RECT  1.995 0.550 2.085 0.810 ;
        RECT  1.825 2.900 2.085 3.160 ;
        RECT  1.835 0.550 1.995 1.425 ;
        RECT  1.825 0.550 1.835 1.045 ;
        RECT  1.225 0.885 1.825 1.045 ;
        RECT  1.775 2.900 1.825 3.080 ;
        RECT  1.615 1.605 1.775 3.080 ;
        RECT  1.565 1.605 1.615 1.765 ;
        RECT  0.895 2.920 1.615 3.080 ;
        RECT  1.405 1.225 1.565 1.765 ;
        RECT  0.885 0.460 1.505 0.620 ;
        RECT  1.275 2.180 1.435 2.600 ;
        RECT  1.225 2.180 1.275 2.340 ;
        RECT  1.065 0.885 1.225 2.340 ;
        RECT  0.885 2.580 1.035 2.740 ;
        RECT  0.635 2.920 0.895 3.180 ;
        RECT  0.725 0.460 0.885 2.740 ;
        RECT  0.615 2.145 0.725 2.405 ;
    END
END TBUFX4

MACRO TBUFX3
    CLASS CORE ;
    FOREIGN TBUFX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  3.045 1.105 3.095 2.585 ;
        RECT  2.885 0.640 3.045 2.860 ;
        RECT  2.785 0.640 2.885 0.900 ;
        RECT  2.785 2.260 2.885 2.860 ;
        END
        ANTENNADIFFAREA     0.6042 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.595 0.505 1.855 ;
        RECT  0.125 1.595 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1118 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.905 2.255 2.400 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 -0.250 3.680 0.250 ;
        RECT  3.295 -0.250 3.555 0.900 ;
        RECT  2.535 -0.250 3.295 0.250 ;
        RECT  2.275 -0.250 2.535 0.900 ;
        RECT  0.385 -0.250 2.275 0.250 ;
        RECT  0.125 -0.250 0.385 0.845 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 3.440 3.680 3.940 ;
        RECT  3.295 2.260 3.555 3.940 ;
        RECT  2.505 3.440 3.295 3.940 ;
        RECT  2.245 2.580 2.505 3.940 ;
        RECT  0.385 3.440 2.245 3.940 ;
        RECT  0.125 2.750 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.070 1.225 2.705 1.385 ;
        RECT  2.655 1.655 2.705 1.915 ;
        RECT  2.445 1.565 2.655 1.915 ;
        RECT  1.775 1.565 2.445 1.725 ;
        RECT  1.910 0.475 2.070 1.385 ;
        RECT  1.775 2.955 1.995 3.215 ;
        RECT  1.215 0.475 1.910 0.735 ;
        RECT  1.615 1.565 1.775 3.215 ;
        RECT  1.575 1.565 1.615 1.725 ;
        RECT  0.715 2.955 1.615 3.215 ;
        RECT  1.415 1.065 1.575 1.725 ;
        RECT  1.275 2.180 1.435 2.600 ;
        RECT  1.215 2.180 1.275 2.340 ;
        RECT  1.055 0.475 1.215 2.340 ;
        RECT  0.875 2.615 1.085 2.775 ;
        RECT  0.715 0.815 0.875 2.775 ;
        RECT  0.690 1.205 0.715 1.485 ;
        RECT  0.615 2.145 0.715 2.405 ;
    END
END TBUFX3

MACRO TBUFX2
    CLASS CORE ;
    FOREIGN TBUFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 0.675 3.095 3.065 ;
        RECT  2.835 0.675 2.885 1.275 ;
        RECT  2.835 2.125 2.885 3.065 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.595 0.460 1.855 ;
        RECT  0.125 1.400 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1001 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.105 2.635 2.175 ;
        RECT  2.425 0.915 2.585 2.545 ;
        RECT  2.065 0.915 2.425 1.075 ;
        RECT  2.115 2.375 2.425 2.545 ;
        RECT  1.955 2.375 2.115 2.635 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 -0.250 3.220 0.250 ;
        RECT  2.295 -0.250 2.555 0.700 ;
        RECT  0.385 -0.250 2.295 0.250 ;
        RECT  0.125 -0.250 0.385 0.855 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 3.440 3.220 3.940 ;
        RECT  2.295 2.725 2.555 3.940 ;
        RECT  0.385 3.440 2.295 3.940 ;
        RECT  0.125 2.750 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.075 1.255 2.235 2.195 ;
        RECT  1.775 1.255 2.075 1.415 ;
        RECT  1.775 2.035 2.075 2.195 ;
        RECT  1.330 0.475 1.885 0.735 ;
        RECT  1.430 1.675 1.805 1.835 ;
        RECT  1.515 1.065 1.775 1.415 ;
        RECT  1.615 2.035 1.775 3.215 ;
        RECT  0.835 2.955 1.615 3.215 ;
        RECT  1.330 1.675 1.430 2.405 ;
        RECT  1.170 0.475 1.330 2.405 ;
        RECT  0.875 2.615 1.115 2.775 ;
        RECT  0.900 0.815 0.955 1.075 ;
        RECT  0.875 0.815 0.900 1.445 ;
        RECT  0.715 0.815 0.875 2.775 ;
        RECT  0.695 0.815 0.715 1.445 ;
        RECT  0.615 2.145 0.715 2.405 ;
        RECT  0.640 1.185 0.695 1.445 ;
    END
END TBUFX2

MACRO TBUFX1
    CLASS CORE ;
    FOREIGN TBUFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.035 3.100 3.060 ;
        RECT  2.835 1.035 2.885 1.295 ;
        RECT  2.835 2.460 2.885 3.060 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 1.545 0.645 1.805 ;
        RECT  0.335 1.645 0.385 1.805 ;
        RECT  0.125 1.645 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0988 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.605 1.695 1.775 2.475 ;
        RECT  1.505 1.695 1.605 2.005 ;
        END
        ANTENNAGATEAREA     0.0468 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 -0.250 3.220 0.250 ;
        RECT  2.285 -0.250 2.545 0.835 ;
        RECT  0.725 -0.250 2.285 0.250 ;
        RECT  0.385 -0.250 0.725 0.405 ;
        RECT  0.125 -0.250 0.385 1.135 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 3.440 3.220 3.940 ;
        RECT  2.325 2.460 2.585 3.940 ;
        RECT  1.985 3.440 2.325 3.940 ;
        RECT  1.725 3.285 1.985 3.940 ;
        RECT  0.385 3.440 1.725 3.940 ;
        RECT  0.125 2.795 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.115 2.020 2.705 2.280 ;
        RECT  2.560 1.410 2.655 1.670 ;
        RECT  2.400 1.015 2.560 1.670 ;
        RECT  2.060 1.015 2.400 1.175 ;
        RECT  2.395 1.410 2.400 1.670 ;
        RECT  1.955 1.355 2.115 2.815 ;
        RECT  1.900 0.870 2.060 1.175 ;
        RECT  1.705 1.355 1.955 1.515 ;
        RECT  1.515 2.655 1.955 2.815 ;
        RECT  1.605 0.870 1.900 1.030 ;
        RECT  1.545 1.225 1.705 1.515 ;
        RECT  1.355 0.655 1.605 1.030 ;
        RECT  1.355 2.655 1.515 3.215 ;
        RECT  1.325 2.195 1.425 2.355 ;
        RECT  1.345 0.655 1.355 1.480 ;
        RECT  0.755 2.955 1.355 3.215 ;
        RECT  1.325 0.870 1.345 1.480 ;
        RECT  1.195 0.870 1.325 2.355 ;
        RECT  1.165 1.320 1.195 2.355 ;
        RECT  0.985 2.565 1.090 2.725 ;
        RECT  0.985 0.695 1.015 0.955 ;
        RECT  0.825 0.695 0.985 2.725 ;
        RECT  0.615 2.145 0.825 2.405 ;
    END
END TBUFX1

MACRO TBUFXL
    CLASS CORE ;
    FOREIGN TBUFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 0.470 2.635 2.820 ;
        RECT  2.425 0.470 2.475 0.760 ;
        RECT  2.375 2.560 2.475 2.820 ;
        RECT  2.375 0.495 2.425 0.755 ;
        END
        ANTENNADIFFAREA     0.2161 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.625 0.505 1.885 ;
        RECT  0.125 1.485 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.785 1.850 2.400 ;
        END
        ANTENNAGATEAREA     0.0468 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.060 -0.250 2.760 0.250 ;
        RECT  1.800 -0.250 2.060 0.405 ;
        RECT  0.385 -0.250 1.800 0.250 ;
        RECT  0.125 -0.250 0.385 0.830 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.010 3.440 2.760 3.940 ;
        RECT  1.750 3.285 2.010 3.940 ;
        RECT  0.385 3.440 1.750 3.940 ;
        RECT  0.125 2.790 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.195 0.940 2.295 1.215 ;
        RECT  2.190 2.120 2.295 2.380 ;
        RECT  2.035 0.800 2.195 1.215 ;
        RECT  2.030 1.395 2.190 3.100 ;
        RECT  1.490 0.800 2.035 0.960 ;
        RECT  1.580 1.395 2.030 1.555 ;
        RECT  1.310 2.940 2.030 3.100 ;
        RECT  1.420 1.235 1.580 1.555 ;
        RECT  1.240 0.605 1.490 0.960 ;
        RECT  0.710 2.940 1.310 3.200 ;
        RECT  1.240 2.155 1.275 2.415 ;
        RECT  1.230 0.605 1.240 2.415 ;
        RECT  1.080 0.800 1.230 2.415 ;
        RECT  0.845 2.600 1.065 2.760 ;
        RECT  0.895 0.430 0.925 0.590 ;
        RECT  0.845 0.430 0.895 1.445 ;
        RECT  0.735 0.430 0.845 2.760 ;
        RECT  0.665 0.430 0.735 0.590 ;
        RECT  0.685 1.185 0.735 2.760 ;
        RECT  0.635 1.185 0.685 1.445 ;
        RECT  0.555 2.155 0.685 2.415 ;
    END
END TBUFXL

MACRO INVX20
    CLASS CORE ;
    FOREIGN INVX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.980 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.715 0.680 4.975 2.980 ;
        RECT  4.490 0.870 4.715 2.775 ;
        RECT  4.015 0.865 4.490 2.775 ;
        RECT  3.955 0.865 4.015 2.995 ;
        RECT  3.805 0.680 3.955 3.150 ;
        RECT  3.695 0.680 3.805 1.280 ;
        RECT  3.695 2.210 3.805 3.150 ;
        RECT  2.935 0.865 3.695 1.280 ;
        RECT  2.935 2.210 3.695 2.775 ;
        RECT  2.675 0.680 2.935 1.280 ;
        RECT  2.675 2.210 2.935 3.150 ;
        RECT  1.915 0.865 2.675 1.280 ;
        RECT  1.915 2.210 2.675 2.775 ;
        RECT  1.655 0.680 1.915 1.280 ;
        RECT  1.655 2.210 1.915 3.150 ;
        RECT  0.895 0.865 1.655 1.280 ;
        RECT  0.895 2.210 1.655 2.775 ;
        RECT  0.635 0.680 0.895 1.280 ;
        RECT  0.635 2.210 0.895 2.810 ;
        RECT  0.585 2.335 0.635 2.585 ;
        END
        ANTENNADIFFAREA     3.9928 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.500 3.585 1.760 ;
        RECT  1.045 1.500 1.255 1.990 ;
        RECT  0.265 1.500 1.045 1.760 ;
        END
        ANTENNAGATEAREA     2.7040 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.490 -0.250 5.980 0.250 ;
        RECT  5.230 -0.250 5.490 1.275 ;
        RECT  4.465 -0.250 5.230 0.250 ;
        RECT  4.205 -0.250 4.465 0.685 ;
        RECT  3.445 -0.250 4.205 0.250 ;
        RECT  3.185 -0.250 3.445 0.685 ;
        RECT  2.425 -0.250 3.185 0.250 ;
        RECT  2.165 -0.250 2.425 0.685 ;
        RECT  1.405 -0.250 2.165 0.250 ;
        RECT  1.145 -0.250 1.405 0.685 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.275 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.490 3.440 5.980 3.940 ;
        RECT  5.230 2.075 5.490 3.940 ;
        RECT  4.465 3.440 5.230 3.940 ;
        RECT  4.205 2.955 4.465 3.940 ;
        RECT  3.445 3.440 4.205 3.940 ;
        RECT  3.185 2.955 3.445 3.940 ;
        RECT  2.425 3.440 3.185 3.940 ;
        RECT  2.165 2.955 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.955 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.075 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END INVX20

MACRO INVX16
    CLASS CORE ;
    FOREIGN INVX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.955 1.105 4.015 2.995 ;
        RECT  3.695 0.680 3.955 3.150 ;
        RECT  2.935 0.865 3.695 2.775 ;
        RECT  2.885 0.680 2.935 3.150 ;
        RECT  2.675 0.680 2.885 1.280 ;
        RECT  2.675 2.210 2.885 3.150 ;
        RECT  1.915 0.865 2.675 1.280 ;
        RECT  1.915 2.210 2.675 2.775 ;
        RECT  1.655 0.680 1.915 1.280 ;
        RECT  1.655 2.210 1.915 3.150 ;
        RECT  0.895 0.865 1.655 1.280 ;
        RECT  0.895 2.210 1.655 2.775 ;
        RECT  0.635 0.680 0.895 1.280 ;
        RECT  0.635 2.210 0.895 2.810 ;
        RECT  0.585 2.335 0.635 2.585 ;
        END
        ANTENNADIFFAREA     3.2232 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.500 2.595 1.760 ;
        RECT  1.045 1.500 1.255 1.990 ;
        RECT  0.295 1.500 1.045 1.760 ;
        END
        ANTENNAGATEAREA     2.1944 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 -0.250 4.600 0.250 ;
        RECT  4.205 -0.250 4.465 1.075 ;
        RECT  3.445 -0.250 4.205 0.250 ;
        RECT  3.185 -0.250 3.445 0.685 ;
        RECT  2.425 -0.250 3.185 0.250 ;
        RECT  2.165 -0.250 2.425 0.685 ;
        RECT  1.405 -0.250 2.165 0.250 ;
        RECT  1.145 -0.250 1.405 0.685 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.275 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 3.440 4.600 3.940 ;
        RECT  4.205 2.275 4.465 3.940 ;
        RECT  3.445 3.440 4.205 3.940 ;
        RECT  3.185 2.955 3.445 3.940 ;
        RECT  2.425 3.440 3.185 3.940 ;
        RECT  2.165 2.955 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.955 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.075 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END INVX16

MACRO INVX12
    CLASS CORE ;
    FOREIGN INVX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 0.680 2.995 2.775 ;
        RECT  2.735 0.680 2.935 3.150 ;
        RECT  2.675 0.915 2.735 3.150 ;
        RECT  2.045 0.915 2.675 2.775 ;
        RECT  1.915 0.680 2.045 2.775 ;
        RECT  1.655 0.680 1.915 3.125 ;
        RECT  1.615 0.680 1.655 2.775 ;
        RECT  0.635 0.680 1.615 1.280 ;
        RECT  0.635 2.175 1.615 2.775 ;
        RECT  0.585 2.335 0.635 2.585 ;
        END
        ANTENNADIFFAREA     2.3948 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.585 1.405 1.845 ;
        RECT  1.045 1.585 1.255 1.990 ;
        RECT  0.465 1.585 1.045 1.845 ;
        END
        ANTENNAGATEAREA     1.6276 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.505 -0.250 3.680 0.250 ;
        RECT  3.245 -0.250 3.505 1.075 ;
        RECT  2.485 -0.250 3.245 0.250 ;
        RECT  2.225 -0.250 2.485 0.735 ;
        RECT  1.435 -0.250 2.225 0.250 ;
        RECT  1.175 -0.250 1.435 0.405 ;
        RECT  0.385 -0.250 1.175 0.250 ;
        RECT  0.125 -0.250 0.385 1.275 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.445 3.440 3.680 3.940 ;
        RECT  3.185 2.275 3.445 3.940 ;
        RECT  2.425 3.440 3.185 3.940 ;
        RECT  2.165 2.955 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.955 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.075 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END INVX12

MACRO INVX8
    CLASS CORE ;
    FOREIGN INVX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.060 0.995 2.635 2.400 ;
        RECT  2.020 0.635 2.060 2.400 ;
        RECT  1.965 0.635 2.020 2.950 ;
        RECT  1.760 0.635 1.965 1.295 ;
        RECT  1.695 1.995 1.965 2.950 ;
        RECT  1.690 0.880 1.760 1.295 ;
        RECT  0.915 1.995 1.695 2.400 ;
        RECT  1.070 0.895 1.690 1.295 ;
        RECT  0.980 0.880 1.070 1.295 ;
        RECT  0.680 0.645 0.980 1.295 ;
        RECT  0.615 1.995 0.915 2.950 ;
        RECT  0.585 2.335 0.615 2.585 ;
        END
        ANTENNADIFFAREA     1.6294 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.515 1.405 1.775 ;
        RECT  0.335 1.615 0.465 1.775 ;
        RECT  0.125 1.615 0.335 1.990 ;
        END
        ANTENNAGATEAREA     1.0868 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 -0.250 2.760 0.250 ;
        RECT  2.325 -0.250 2.585 0.745 ;
        RECT  1.500 -0.250 2.325 0.250 ;
        RECT  1.240 -0.250 1.500 0.405 ;
        RECT  0.420 -0.250 1.240 0.250 ;
        RECT  0.160 -0.250 0.420 1.185 ;
        RECT  0.000 -0.250 0.160 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 3.440 2.760 3.940 ;
        RECT  2.285 2.755 2.545 3.940 ;
        RECT  1.435 3.440 2.285 3.940 ;
        RECT  1.175 2.615 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END INVX8

MACRO INVX6
    CLASS CORE ;
    FOREIGN INVX6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.060 1.105 2.175 2.585 ;
        RECT  1.725 0.670 2.060 2.900 ;
        RECT  1.700 0.980 1.725 2.900 ;
        RECT  1.045 0.980 1.700 2.375 ;
        RECT  0.945 0.980 1.045 1.280 ;
        RECT  0.945 2.075 1.045 2.375 ;
        RECT  0.645 0.625 0.945 1.280 ;
        RECT  0.645 2.075 0.945 3.185 ;
        RECT  0.585 2.335 0.645 2.995 ;
        END
        ANTENNADIFFAREA     1.5283 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.495 1.545 0.755 1.805 ;
        RECT  0.335 1.545 0.495 1.705 ;
        RECT  0.175 1.290 0.335 1.705 ;
        RECT  0.125 1.290 0.175 1.580 ;
        END
        ANTENNAGATEAREA     0.8268 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 -0.250 2.300 0.250 ;
        RECT  1.205 -0.250 1.465 0.800 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 1.090 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 3.440 2.300 3.940 ;
        RECT  1.205 2.555 1.465 3.940 ;
        RECT  0.385 3.440 1.205 3.940 ;
        RECT  0.125 2.200 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END INVX6

MACRO INVX4
    CLASS CORE ;
    FOREIGN INVX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.025 1.290 1.255 1.990 ;
        RECT  0.765 0.695 1.025 2.915 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.450 0.555 1.830 ;
        RECT  0.135 1.450 0.335 1.990 ;
        RECT  0.125 1.700 0.135 1.990 ;
        END
        ANTENNAGATEAREA     0.5512 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 -0.250 1.840 0.250 ;
        RECT  1.305 -0.250 1.565 1.110 ;
        RECT  0.485 -0.250 1.305 0.250 ;
        RECT  0.225 -0.250 0.485 1.200 ;
        RECT  0.000 -0.250 0.225 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 3.440 1.840 3.940 ;
        RECT  1.305 2.210 1.565 3.940 ;
        RECT  0.485 3.440 1.305 3.940 ;
        RECT  0.225 2.195 0.485 3.940 ;
        RECT  0.000 3.440 0.225 3.940 ;
        END
    END VDD
END INVX4

MACRO INVX3
    CLASS CORE ;
    FOREIGN INVX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.380 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.205 1.355 1.255 2.175 ;
        RECT  1.045 1.285 1.205 2.330 ;
        RECT  0.795 1.285 1.045 1.445 ;
        RECT  0.795 2.170 1.045 2.330 ;
        RECT  0.785 1.105 0.795 1.445 ;
        RECT  0.785 2.170 0.795 2.585 ;
        RECT  0.625 0.980 0.785 1.445 ;
        RECT  0.525 2.170 0.785 2.770 ;
        RECT  0.525 0.980 0.625 1.240 ;
        END
        ANTENNADIFFAREA     0.5776 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.530 1.625 0.790 1.885 ;
        RECT  0.335 1.700 0.530 1.885 ;
        RECT  0.125 1.700 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.3952 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 -0.250 1.380 0.250 ;
        RECT  0.995 -0.250 1.255 0.405 ;
        RECT  0.385 -0.250 0.995 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 3.440 1.380 3.940 ;
        RECT  0.995 3.285 1.255 3.940 ;
        RECT  0.385 3.440 0.995 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END INVX3

MACRO INVX2
    CLASS CORE ;
    FOREIGN INVX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.380 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 1.105 1.255 2.585 ;
        RECT  0.920 0.595 1.080 3.115 ;
        RECT  0.820 0.595 0.920 1.295 ;
        RECT  0.820 2.175 0.920 3.115 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.585 0.735 1.990 ;
        RECT  0.125 1.700 0.475 1.990 ;
        END
        ANTENNAGATEAREA     0.2756 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 -0.250 1.380 0.250 ;
        RECT  0.280 -0.250 0.540 1.225 ;
        RECT  0.000 -0.250 0.280 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 3.440 1.380 3.940 ;
        RECT  0.280 2.215 0.540 3.940 ;
        RECT  0.000 3.440 0.280 3.940 ;
        END
    END VDD
END INVX2

MACRO INVX1
    CLASS CORE ;
    FOREIGN INVX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 1.105 0.795 2.585 ;
        RECT  0.585 1.035 0.785 2.715 ;
        RECT  0.525 1.035 0.585 1.295 ;
        RECT  0.525 2.115 0.585 2.715 ;
        END
        ANTENNADIFFAREA     0.3604 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.515 0.405 1.935 ;
        RECT  0.125 1.515 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.250 0.920 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 0.920 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END INVX1

MACRO INVXL
    CLASS CORE ;
    FOREIGN INVXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 1.290 0.795 2.400 ;
        RECT  0.745 1.290 0.785 2.510 ;
        RECT  0.585 1.035 0.745 2.510 ;
        RECT  0.385 1.035 0.585 1.295 ;
        RECT  0.525 2.250 0.585 2.510 ;
        END
        ANTENNADIFFAREA     0.2265 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.555 0.405 2.065 ;
        END
        ANTENNAGATEAREA     0.0728 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.605 -0.250 0.920 0.250 ;
        RECT  0.345 -0.250 0.605 0.405 ;
        RECT  0.000 -0.250 0.345 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 0.920 3.940 ;
        RECT  0.125 2.875 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END INVXL

MACRO BUFX20
    CLASS CORE ;
    FOREIGN BUFX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.015 0.695 7.135 2.010 ;
        RECT  6.875 0.695 7.015 3.005 ;
        RECT  6.755 1.020 6.875 3.005 ;
        RECT  6.115 1.020 6.755 2.400 ;
        RECT  5.995 0.585 6.115 2.400 ;
        RECT  5.855 0.585 5.995 3.115 ;
        RECT  5.735 1.020 5.855 3.115 ;
        RECT  5.165 1.020 5.735 2.400 ;
        RECT  4.975 0.585 5.165 2.400 ;
        RECT  4.715 0.585 4.975 2.895 ;
        RECT  4.525 0.585 4.715 2.435 ;
        RECT  2.675 0.585 4.525 1.185 ;
        RECT  3.955 1.845 4.525 2.435 ;
        RECT  3.695 1.845 3.955 2.895 ;
        RECT  2.935 1.845 3.695 2.435 ;
        RECT  2.675 1.845 2.935 2.895 ;
        END
        ANTENNADIFFAREA     4.0075 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.645 1.405 1.905 ;
        RECT  0.335 1.700 0.465 1.905 ;
        RECT  0.125 1.700 0.335 1.990 ;
        END
        ANTENNAGATEAREA     1.0634 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.645 -0.250 7.820 0.250 ;
        RECT  7.385 -0.250 7.645 1.275 ;
        RECT  6.625 -0.250 7.385 0.250 ;
        RECT  6.365 -0.250 6.625 0.755 ;
        RECT  5.605 -0.250 6.365 0.250 ;
        RECT  5.345 -0.250 5.605 0.755 ;
        RECT  4.555 -0.250 5.345 0.250 ;
        RECT  4.295 -0.250 4.555 0.405 ;
        RECT  3.475 -0.250 4.295 0.250 ;
        RECT  3.215 -0.250 3.475 0.405 ;
        RECT  2.425 -0.250 3.215 0.250 ;
        RECT  2.165 -0.250 2.425 1.125 ;
        RECT  1.405 -0.250 2.165 0.250 ;
        RECT  1.145 -0.250 1.405 1.125 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.125 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.525 3.440 7.820 3.940 ;
        RECT  7.265 2.405 7.525 3.940 ;
        RECT  6.505 3.440 7.265 3.940 ;
        RECT  6.245 2.615 6.505 3.940 ;
        RECT  5.485 3.440 6.245 3.940 ;
        RECT  5.225 2.615 5.485 3.940 ;
        RECT  4.465 3.440 5.225 3.940 ;
        RECT  4.205 2.615 4.465 3.940 ;
        RECT  3.445 3.440 4.205 3.940 ;
        RECT  3.185 2.615 3.445 3.940 ;
        RECT  2.425 3.440 3.185 3.940 ;
        RECT  2.165 2.275 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.615 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.915 1.455 4.125 1.615 ;
        RECT  1.755 0.695 1.915 3.120 ;
        RECT  1.655 0.695 1.755 1.465 ;
        RECT  1.655 2.180 1.755 3.120 ;
        RECT  0.895 1.305 1.655 1.465 ;
        RECT  0.895 2.180 1.655 2.340 ;
        RECT  0.735 0.695 0.895 1.465 ;
        RECT  0.635 2.180 0.895 3.120 ;
        RECT  0.635 0.695 0.735 1.295 ;
    END
END BUFX20

MACRO BUFX16
    CLASS CORE ;
    FOREIGN BUFX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.650 1.290 6.315 2.400 ;
        RECT  5.470 0.655 5.650 2.400 ;
        RECT  5.210 0.655 5.470 2.720 ;
        RECT  5.185 0.655 5.210 2.585 ;
        RECT  4.965 0.655 5.185 2.455 ;
        RECT  2.165 0.655 4.965 1.255 ;
        RECT  4.475 1.855 4.965 2.455 ;
        RECT  4.465 1.855 4.475 2.585 ;
        RECT  4.205 1.855 4.465 2.895 ;
        RECT  3.445 1.855 4.205 2.455 ;
        RECT  3.185 1.855 3.445 2.895 ;
        RECT  2.425 1.855 3.185 2.455 ;
        RECT  2.165 1.855 2.425 2.895 ;
        END
        ANTENNADIFFAREA     3.0144 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.580 1.510 1.840 ;
        RECT  0.585 1.580 0.795 1.990 ;
        RECT  0.570 1.580 0.585 1.840 ;
        END
        ANTENNAGATEAREA     0.8424 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.130 -0.250 6.440 0.250 ;
        RECT  5.870 -0.250 6.130 1.065 ;
        RECT  5.125 -0.250 5.870 0.250 ;
        RECT  4.865 -0.250 5.125 0.405 ;
        RECT  4.045 -0.250 4.865 0.250 ;
        RECT  3.785 -0.250 4.045 0.405 ;
        RECT  2.965 -0.250 3.785 0.250 ;
        RECT  2.705 -0.250 2.965 0.405 ;
        RECT  1.915 -0.250 2.705 0.250 ;
        RECT  1.655 -0.250 1.915 0.955 ;
        RECT  0.895 -0.250 1.655 0.250 ;
        RECT  0.635 -0.250 0.895 0.935 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.010 3.440 6.440 3.940 ;
        RECT  5.750 2.895 6.010 3.940 ;
        RECT  5.005 3.440 5.750 3.940 ;
        RECT  4.745 3.285 5.005 3.940 ;
        RECT  3.955 3.440 4.745 3.940 ;
        RECT  3.695 2.635 3.955 3.940 ;
        RECT  2.935 3.440 3.695 3.940 ;
        RECT  2.675 2.635 2.935 3.940 ;
        RECT  1.915 3.440 2.675 3.940 ;
        RECT  1.655 2.610 1.915 3.940 ;
        RECT  0.895 3.440 1.655 3.940 ;
        RECT  0.635 2.605 0.895 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.945 1.475 4.745 1.635 ;
        RECT  1.785 1.240 1.945 2.400 ;
        RECT  1.405 1.240 1.785 1.400 ;
        RECT  1.405 2.240 1.785 2.400 ;
        RECT  1.145 0.695 1.405 1.400 ;
        RECT  1.145 2.240 1.405 3.180 ;
        RECT  0.385 1.240 1.145 1.400 ;
        RECT  0.385 2.240 1.145 2.400 ;
        RECT  0.125 0.695 0.385 1.400 ;
        RECT  0.125 2.240 0.385 3.180 ;
    END
END BUFX16

MACRO BUFX12
    CLASS CORE ;
    FOREIGN BUFX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.955 1.105 4.015 2.585 ;
        RECT  3.695 0.880 3.955 2.875 ;
        RECT  3.305 0.880 3.695 2.640 ;
        RECT  2.935 0.880 3.305 1.385 ;
        RECT  2.935 2.040 3.305 2.640 ;
        RECT  2.675 0.645 2.935 1.385 ;
        RECT  2.675 2.040 2.935 3.045 ;
        RECT  1.915 0.880 2.675 1.385 ;
        RECT  1.915 2.040 2.675 2.640 ;
        RECT  1.655 0.645 1.915 1.385 ;
        RECT  1.655 2.040 1.915 3.045 ;
        END
        ANTENNADIFFAREA     2.4024 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.595 1.065 1.755 ;
        RECT  0.150 1.595 0.335 1.990 ;
        RECT  0.125 1.700 0.150 1.990 ;
        END
        ANTENNAGATEAREA     0.5616 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 -0.250 4.600 0.250 ;
        RECT  4.205 -0.250 4.465 1.275 ;
        RECT  3.445 -0.250 4.205 0.250 ;
        RECT  3.185 -0.250 3.445 0.685 ;
        RECT  2.425 -0.250 3.185 0.250 ;
        RECT  2.165 -0.250 2.425 0.685 ;
        RECT  1.405 -0.250 2.165 0.250 ;
        RECT  1.145 -0.250 1.405 1.075 ;
        RECT  0.385 -0.250 1.145 0.250 ;
        RECT  0.125 -0.250 0.385 1.075 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 3.440 4.600 3.940 ;
        RECT  4.205 2.075 4.465 3.940 ;
        RECT  3.445 3.440 4.205 3.940 ;
        RECT  3.185 2.955 3.445 3.940 ;
        RECT  2.425 3.440 3.185 3.940 ;
        RECT  2.165 2.955 2.425 3.940 ;
        RECT  1.405 3.440 2.165 3.940 ;
        RECT  1.145 2.275 1.405 3.940 ;
        RECT  0.385 3.440 1.145 3.940 ;
        RECT  0.125 2.275 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.420 1.605 3.105 1.765 ;
        RECT  1.260 1.255 1.420 2.095 ;
        RECT  0.895 1.255 1.260 1.415 ;
        RECT  0.895 1.935 1.260 2.095 ;
        RECT  0.635 0.695 0.895 1.415 ;
        RECT  0.635 1.935 0.895 2.910 ;
    END
END BUFX12

MACRO BUFX8
    CLASS CORE ;
    FOREIGN BUFX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.025 1.105 3.095 2.585 ;
        RECT  2.765 0.695 3.025 2.895 ;
        RECT  2.425 1.020 2.765 2.475 ;
        RECT  1.945 1.020 2.425 1.355 ;
        RECT  1.945 1.995 2.425 2.475 ;
        RECT  1.685 0.695 1.945 1.355 ;
        RECT  1.685 1.995 1.945 2.935 ;
        END
        ANTENNADIFFAREA     1.6112 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.615 1.010 1.775 ;
        RECT  0.125 1.615 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.4212 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.535 -0.250 3.680 0.250 ;
        RECT  3.275 -0.250 3.535 1.095 ;
        RECT  2.485 -0.250 3.275 0.250 ;
        RECT  2.225 -0.250 2.485 0.795 ;
        RECT  1.435 -0.250 2.225 0.250 ;
        RECT  1.175 -0.250 1.435 1.095 ;
        RECT  0.385 -0.250 1.175 0.250 ;
        RECT  0.125 -0.250 0.385 1.295 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.535 3.440 3.680 3.940 ;
        RECT  3.275 2.255 3.535 3.940 ;
        RECT  2.485 3.440 3.275 3.940 ;
        RECT  2.225 2.875 2.485 3.940 ;
        RECT  1.435 3.440 2.225 3.940 ;
        RECT  1.175 2.295 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.295 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.475 1.545 2.115 1.805 ;
        RECT  1.315 1.275 1.475 2.115 ;
        RECT  0.895 1.275 1.315 1.435 ;
        RECT  0.895 1.955 1.315 2.115 ;
        RECT  0.635 0.695 0.895 1.435 ;
        RECT  0.635 1.955 0.895 2.555 ;
    END
END BUFX8

MACRO BUFX6
    CLASS CORE ;
    FOREIGN BUFX6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.025 2.335 3.095 2.585 ;
        RECT  2.765 0.675 3.025 1.275 ;
        RECT  2.765 1.975 3.025 2.915 ;
        RECT  2.635 0.975 2.765 1.275 ;
        RECT  2.635 1.975 2.765 2.345 ;
        RECT  1.965 0.975 2.635 2.345 ;
        RECT  1.945 0.975 1.965 1.275 ;
        RECT  1.945 1.975 1.965 2.345 ;
        RECT  1.685 0.675 1.945 1.275 ;
        RECT  1.685 1.975 1.945 2.915 ;
        END
        ANTENNADIFFAREA     1.5280 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.595 1.055 1.755 ;
        RECT  0.125 1.595 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.3198 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 -0.250 3.220 0.250 ;
        RECT  2.225 -0.250 2.485 0.795 ;
        RECT  1.435 -0.250 2.225 0.250 ;
        RECT  1.175 -0.250 1.435 1.075 ;
        RECT  0.385 -0.250 1.175 0.250 ;
        RECT  0.125 -0.250 0.385 1.085 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 3.440 3.220 3.940 ;
        RECT  2.225 2.555 2.485 3.940 ;
        RECT  1.435 3.440 2.225 3.940 ;
        RECT  1.175 2.420 1.435 3.940 ;
        RECT  0.385 3.440 1.175 3.940 ;
        RECT  0.125 2.170 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.470 1.510 1.775 1.770 ;
        RECT  1.310 1.255 1.470 2.100 ;
        RECT  0.895 1.255 1.310 1.415 ;
        RECT  0.895 1.940 1.310 2.100 ;
        RECT  0.635 1.010 0.895 1.415 ;
        RECT  0.635 1.940 0.895 2.670 ;
    END
END BUFX6

MACRO BUFX4
    CLASS CORE ;
    FOREIGN BUFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.160 1.290 2.175 1.990 ;
        RECT  2.155 1.095 2.160 1.990 ;
        RECT  1.960 1.095 2.155 2.170 ;
        RECT  1.535 1.095 1.960 1.295 ;
        RECT  1.955 1.540 1.960 2.170 ;
        RECT  1.690 1.970 1.955 2.170 ;
        RECT  1.575 1.970 1.690 2.175 ;
        RECT  1.315 1.970 1.575 2.910 ;
        RECT  1.275 0.695 1.535 1.295 ;
        END
        ANTENNADIFFAREA     0.8904 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.795 1.770 ;
        RECT  0.485 1.510 0.585 1.770 ;
        END
        ANTENNAGATEAREA     0.2132 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 -0.250 2.300 0.250 ;
        RECT  1.855 -0.250 2.115 0.795 ;
        RECT  0.995 -0.250 1.855 0.250 ;
        RECT  0.735 -0.250 0.995 1.085 ;
        RECT  0.000 -0.250 0.735 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 3.440 2.300 3.940 ;
        RECT  1.855 2.555 2.115 3.940 ;
        RECT  0.995 3.440 1.855 3.940 ;
        RECT  0.735 2.305 0.995 3.940 ;
        RECT  0.000 3.440 0.735 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.135 1.510 1.705 1.770 ;
        RECT  0.975 1.510 1.135 2.115 ;
        RECT  0.405 1.955 0.975 2.115 ;
        RECT  0.305 0.695 0.405 1.295 ;
        RECT  0.305 1.955 0.405 2.895 ;
        RECT  0.145 0.695 0.305 2.895 ;
    END
END BUFX4

MACRO BUFX3
    CLASS CORE ;
    FOREIGN BUFX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 1.135 2.175 1.765 ;
        RECT  1.965 1.135 2.125 2.220 ;
        RECT  1.535 1.135 1.965 1.295 ;
        RECT  1.535 2.060 1.965 2.220 ;
        RECT  1.275 1.035 1.535 1.295 ;
        RECT  1.325 2.060 1.535 2.660 ;
        RECT  1.275 2.400 1.325 2.660 ;
        END
        ANTENNADIFFAREA     0.6042 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.795 1.810 ;
        RECT  0.535 1.550 0.585 1.810 ;
        END
        ANTENNAGATEAREA     0.1612 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.075 -0.250 2.300 0.250 ;
        RECT  1.815 -0.250 2.075 0.795 ;
        RECT  0.995 -0.250 1.815 0.250 ;
        RECT  0.735 -0.250 0.995 1.085 ;
        RECT  0.000 -0.250 0.735 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.075 3.440 2.300 3.940 ;
        RECT  1.815 2.525 2.075 3.940 ;
        RECT  0.995 3.440 1.815 3.940 ;
        RECT  0.735 2.525 0.995 3.940 ;
        RECT  0.000 3.440 0.735 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.135 1.550 1.705 1.810 ;
        RECT  0.975 1.550 1.135 2.200 ;
        RECT  0.455 2.040 0.975 2.200 ;
        RECT  0.355 2.040 0.455 2.640 ;
        RECT  0.355 1.035 0.405 1.295 ;
        RECT  0.195 1.035 0.355 2.640 ;
    END
END BUFX3

MACRO BUFX2
    CLASS CORE ;
    FOREIGN BUFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.665 1.290 1.715 2.175 ;
        RECT  1.505 1.125 1.665 2.370 ;
        RECT  1.315 1.125 1.505 1.285 ;
        RECT  1.315 2.210 1.505 2.370 ;
        RECT  1.055 1.025 1.315 1.285 ;
        RECT  1.055 2.210 1.315 2.470 ;
        END
        ANTENNADIFFAREA     0.4228 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.745 0.880 0.795 1.355 ;
        RECT  0.585 0.880 0.745 1.665 ;
        RECT  0.455 1.405 0.585 1.665 ;
        END
        ANTENNAGATEAREA     0.1053 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 -0.250 1.840 0.250 ;
        RECT  0.635 -0.250 1.715 0.405 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 3.440 1.840 3.940 ;
        RECT  0.795 3.285 1.715 3.940 ;
        RECT  0.000 3.440 0.795 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.215 1.510 1.315 1.770 ;
        RECT  1.055 1.510 1.215 2.030 ;
        RECT  0.385 1.870 1.055 2.030 ;
        RECT  0.275 0.435 0.385 0.695 ;
        RECT  0.275 1.870 0.385 3.050 ;
        RECT  0.115 0.435 0.275 3.050 ;
    END
END BUFX2

END LIBRARY

